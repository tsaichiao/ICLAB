
// `include "../00_TESTBED/pseudo_DRAM.sv"
`include "Usertype.sv"
`define SEEDS 5487
`define PAT_NUM_ 100000


program automatic PATTERN(input clk, INF.PATTERN inf);

`protected
AJ<aQ:&))8<55Q5>D-f]db.><3Z1?6ZSUgbT2VG)=2Q4Q?G;Y8e^4)+V8U1U3J&[
fdXFfM?ReG-7KV_Mg6NC;]ZHT0fPDgSUe2I>52I/+VgFA;#e?R,E5b8gXQCH3bY-
e:A5B>f9aKDD;PgP[HWX13Nc8#[E0QZ.=?N_B>\@G=H&&5Q](PZY#b29d9.gC2D@
NEJI31b+W/aac\/-d\(>c\aac(VG@CLQ5VW=];H_a/UE^^M/<bAIQT+9f>^DP3B-
X;(DZM6H@Ec^@9PF&Z.<E0]EF=ZL^S1Fb_U28-d_g9YIBdG+W367&12cXK^eFJMX
/<-fgCYJW@6d#_ffcb_:T:d\&NIDL(3SbTB?BO+_COdAREQ7cB@83#Tf<\McNYMZ
<E>DN]/\1Ka8+fI1[WgC(K(/-/_0aeR;+LGWYA@@?+S2DOCJCQP?;2O]P^-a3>NN
BgOUbNT<H4+BKO;XAVPTD(Tg(b:&3L-g)6#)R44#<LfR1ZFCLC51Vc3-]6Y?IBWF
D-K-7XLO]AE\HKf:Na7\gJ6OfJ+>KOOG4&D9+7&82I<Z+Z0O5BNCaS[C+A=9aJJ+
ccd<CcffTCc]E<f,#B55;:ZIdbOQ+#fNWC#;ONc:2gc1OZWAL\eYU>E_1PTEU6JM
C36YDXabfUUd8G=FES?H77.UKRGF2g5JF?8-UcS@[:EKJXEGA&HAP<3KZO-d,c@]
&O,=\.+7DX\?f01.,_2)-;<UScL\EHeQAZ9T<[gV1?Q/U/4e&>/SK_\b36QAG#H4
FP4=WY=C5#=7,5[I[MaO<aP=f\3J^J4>U2Y+e2=X[>L_A9R?]GNgBCQE-9VN)a1D
E=A,8CR;cBg(:6P&@2BMEYU?;J6W_C:e7gdM;H3#O>U+[=df4@EV)c90[;B&3Z(C
g^I?g-M1,.Q\5#1cb/Z;D76/0e4Y/6^d_4))1eA^1F5b3:Q(Z?;6PEF]TgWZAMaJ
g=5183Gc//:9X=6Ig(\CZ,QD;C+8B@+95_^W^P#;>J4#ddQ2NHA]>J(>6EB6DM;5
2CT=0=C5-AC:Ka&SZ/71aMMf<A#:R^)?0fX[MVJ-#OT>QD6=C(B)XPYB<PN(M(]X
([Qb<aRdY@PJ_JT&4b[1c4GZ=+Y92eg68]S.V0-][21/G3dO]OIXJ>CQVPb3MQ<8
&OZN9WL.g<3;VW+@L[U6QA)]X&E6\U&g4g?cVPg03(4+@(+e2]Q8eGbC=5\A_J&?
HWY04O\Pe\c:(::?C_:#)d&7Jb8X@I7.gSe)K^SbBGZF->M#J]^BB2dUJE:79faZ
Q;d?N76f-)OECFgOGFI9#W_Z<Wg2>g;(]X_:KZ6\\VY)U@XdcF?.<N#P=M9bK6g2
5CA)CQWK,EVSNG/KDUJ.R9Md/FHMaV52(]V_<ffF7>=IK.g6A5HWVfAT?.H&4E4:
=4D;1Z6ZOb5UZ>,;&A:#1QC>H9&O_M<[IQ0>1S[ge;HQ#N^aKJ32B>WPae0N;A9:
EKUBZgU4S,2=8]8MOOgL6N]1Q2E65c_[TF<L)XE0RAaf5CMV\3IX[]RX.eb9HV;T
ed.=&NZ?CFI^80HR_QBIgK<1(9S<N<gBS(LaT@V0&c=X@C<2)8gM7RK;,^:KN3Z;
4181(>+)C5G^ObA/9C(HMeD>I;9=@A8Y:bK)4V[WFPNWGYZW.=AI#T?\A3M/;.0c
&/@ZS&[MSF>->/GKYZdT\46c[cdI:-[SHCM=(E]X\fPFdB=V2_T8TR=TL^#M,C++
.EU>^3Q1E^?L&<De-1Y7[[CM_B(/VRE4V3A?JMURK([(T,a;Ec6M)?RH_KdMb5YK
HP^g9[[2GfSTESAS+1_IOffZ+aJT-P3f_O-R.c3XfYU0@53#dBB:B@\c1(b/RDcX
Ea/.1RMFB4IL>QM-/+>:Ed=\MeM;/TaKM?O>Ca>M\[(+X;)AL)>B#C[WJfGJcb(9
.&7P98)_]g4)-a-1U#K&KSRONEGWUcP6\9Y+=0gO663#502)1\JHD/KCcVM-cZeX
]/44K\2Q?MX;&M-eN_KQ1a&[H3\JgBYRM<5T&NO)Y:7IL;a7D5?-:Be+0WIScN;g
0g+@&15f&176.58Ka>f>Oed@-?^f(a^5G01(d6#?1).H^O\&YM_5eSgN>P90B(56
,#X/7_LNP\cV=OD9d+VX3Q^aSQ[Q@fTf)A]IX9VG3(YeJE#Vg@?#f&G<G&BN^Z=[
/<SV5F\.N44-DIDb,[WO6\=/5a0Y0R<&WLCeCSN>OPCA#J([gcI,4AC<_5EVP87&
R-6Q[+W9;[13TFYY<gM,f0eG139[>&(IO4D&MSCR^,W9Y2R(b]57)3OQEVHN8LWC
/dA;@.f:df\7YDeb3@U>9^6^B3Q#bKOASUHIcZJgLU@6dG#DBGNH4##ISc?.S<WC
&<<J3)IJ1/OR==98?BN5RLB6111AAJ_M9F>7/Db<REKGB9+)<W7c-#4LUJV,SW_E
Z&PJ1:3U_=5aA+GY=gF>S,B;:@G7C1T+#W9c9D7_PC0P6T^[BQ/aVf2+>2AKP--f
3?d<?5>5gTQaCY)9.3?8QFdPAd=Af_4VWK<[eXYO_cSK4XBQ.8+,gSMgBR/EJeQX
1e)6SAY<WcC\+#aZ(O.-:.5DSL(bM4I;./)fAeE58T.EF4)G/gP[(AS6d/[->7_O
GA.64CccU;+LbXVE=GCbWRWETRVYW)46(HVQb[QGeS5L3A9e]VNP&V_81#->;&RG
/3+G<XE?W#/Q[F0QE>4R4PQK[dZ6#5_9E^HAH6(\IVcH:GJSQ1ILLQ@SPDY>I8GV
[;?<2:+Pc+#JJ+]+0LZ?1,.DD]Q04X)VdPV(Ig0T9OJ3APdZ-3/cMDH?@bXa1aFB
9^UT4MQHC@+SRJD_aQ]8<e^c-1YPa&#Y+6&&1_8MV&7B@AO\,/.]F<U<^@#O?PZc
PN,UOLW@6I1d9RP#^(+AG=LLVc_/H+PPNRbWaH;R@NVXC9d,KA6Q@S07L.]_I8gT
(QHCdB:,9e8I9N:L)Q4gBZZL4QAe=gD9TT8(\Q[Z89DO_DaF/\1YDRLQ\:LF=7Ff
_,?<?+d;(4]8N;aQZY)Me:WTTPSI?f.@b,2GagVGdD;Vf-7((GDb3KPZ0_YMa11S
^b[=gB=,<7R5]-eVC;D994&WS/QO0L=9Z1JK]cbI#aEUL<;C^gS=&#52fQ#DH\Ce
P[3^SR]I?3TL0?@TR3+C>O#\[-Q\2&)=K0C(@4bND05d+_A-B9RZ7@/]^EF^.cdK
f64X^[DgFSbgM.?KWB:F.Dd,DgN\IM7RNQOX(cC8TPQEBK13T\TBQ<+P,XZ3?LCR
Zb>;2R.[H.I3E]Z=8S#WJZ>b-=BJ:TN<6(-Tf\:bT>?Tb;/-gIb_+acCT.#ZE3<_
E.<#dYB>g)MOLB7@-bJ74cb<E0#2,AYH_&2Rb&e<6d=e-[T^CB._;g5C+A.O.;ff
,<a[XB&CLDcF=1.#\G7&RfNRV<(d6ZXAK(Va1TH-8bJ[TKQNMGX<=G)T:AO9=@Kf
._&2?KS5F9V^Qc+1ce@T(LY?79a]6R4Z?BDMa_Z4_923[fV6EO3YZ:YF=6JfaEVE
9IgcYH2&b\+0..@WB\:QZ0:QES2^c_GIGcI#]G(X#RZGL9g;X4KGBF\:Z/4)IWRB
[JWN]f[6RY<@W,cRVJYYN2@@7L?ZD6T2badPbQ9#1#D3\B?/8;7dW/Ke>DUMc(CV
VYb=S^(GL^H)QdN]/-[-VV[8J_P=?>XVMD@4M<e[\B;[(A1;ac7---=b]L4JQ?&G
:?VX2]<M#=Ld_ga]&OV>XWY<FW4Ma3KZL)#aeYCC/U><UU&>;\,K]]8XO.3<-I8V
^R2DXJ,PQMI?BEONSgUWKL;U6V+I:<S^>=a4+A0G/NJS28=X(2>S+@]41YO2GF8O
g71I7)c20M1)8,bd^]KEE_O_U9T(c?&B?AI-f1^;@<B2dbfO1CU4gAf5O2(\ZZ2,
8O^UIHS>2:U6f<L.7K@X^c8=#R6(+a(^S)?3d@1ZPTK_TedL6FZ7W;80K;=SU1TH
K/4K+Gc6]Uf-([<ASW&4N>bBd:=+:\8R1\ED7(C0B+,UQC8]SO>TbC-4X_066&>0
Q>f]A^=:4D)ZVe]TLE,T-82daKeHd=>78f<Y,0VNX<N9A]a]?8N:9aHNE]CX)G0V
TAdHV=2]3cREbc7(g.0?,]FIAc5XcUd]\IG>Kd>Xe5)T9cb,>KF([-??&bLCEI<H
AT/<I<_,CeV=M5b?dFcf+1@[;R+S3NT:I&9I@H#Ae;eORCI18cAI3>cNc\NN;@YQ
T/(^Z.)BI_U/5;ONJa9&a,:L_a<M-??LIgg5E\<aI(M#VGAG=cXV],3JOf:D<<45
48+>#N#Q.G1;ag2Wd2LOe1N5PIZR9S3eBJ.Q+HB.BLZ+f2MS:LWf7^X.MbcWL[#=
LbEG>7P_3V7C2YUT245DQe=<_TT5(]^IM.8F-[d&?N:@SZGP.)\HAX?GNUg_(;F:
^83.H\LT6_I[CMb=W68Zb[>aDO#?V(ED/?bER+;INA>IWR1M-<6VONA3R\ZSN70J
:b(KQH(0MW>0)8NOVXHH=+XF+L]<#@65\O&U-9_KY,gF[a[DPE>3959^?\<6EN=1
O)AP2X6-.2:?=SOU#Z>N_(8-V,V83;-C?A8VN\9H?##fVB+]929\ULAgF7:fcU1]
.eEC\7cL7)59N/Lg?_T5#aM&G)V?AWP(N=+J?S2b38A5A]S/R9.2:RDdAI:+9)g<
S+1,_?,eM?]4YR^[+6[]TdG&D-DY0;E&7UF#GdS\aGLAfYR[[D/3_\d(W5?>V5AH
g&I5(I]gZ^1^Fd265[gRcR[M\gcb)J8^PVggOJ<1]_M:O(#_>b#\EgBO2\)XC]Q1
A>[J-,8]ED00aY#Y#,GBcS;A7@b(JW.O2eX;=8cC6>-P35RG0Lgc.T_fXfPFB:9\
REBKJXVO+>d-V1K@]NB[aXC^Y77/G/E])?[SF;LKBTU?3?7Y1VK:JX90HC2f=RM[
/0;GH#&g5gdMgdCfH\(&9:<AD]b4/fB_VN5,.,4WWfY[C<<DKB26-(Q01I^2E?CH
LTFDSH)Z?26eeG[O;fZb<bf&/,A]/Ga#c;2G)FR#\H5g;>fMA8b0U52S1RI8+BLe
Nb2PTK#>A]KZ3<FC[P@B3#_eNbSLYI8Pe03KW9g7\C2&,6J?:A#DIJM>7SJZ&cK@
A5C0\bH]g5:A#1Z4?4XZT62]4^[fFCLGLO;>\9Rd[a-V@P9,P+VU^HD8bR3>1T_L
YX7e?,_4g(&I74Xf_R#V:^0/N[[cL.7/0ENY_NM/_1>9)1L6F^F61P#R^dM9K6;L
@;_3gF2,H#378:H7KaSB2b/g;g7^aQ=ERANPA0_+[4G\28YRbRUg-:8d^fIfH8Ja
_SEXV<H5-.?UeXUT#6JI0OHWR546:O&0^^218(CafcM&P=R,?W^Q\R\[W_-RE<>:
,.Q9(6MJX+5+]C=NS\XO-8>acU?4dK6d=[PGe&<G7Y,ZPMa/VMHJ]&1c)T2^13+T
TePJHR3X;>(=Ba_XE[Be<Y_DEJM5.J865K1;1Rf2R[OP=#(BQN\27W\d]].L8;7.
#@350>ROTA>^^A^9,=,c6?WdM:_c9cI_6^F5@9=9IR?5Z_a:V_QeA?:4^TJ:G496
X93@Z@Cf60P9cWKH[&dO]9VcGK]5V<N390A?E9POJL\8:WCSBa5K\W)Pd5Jcc5>T
M[W8N(CeFM)U6E]KaEFJU4QFgX\K<DBNGF?)TF)-:aB<[M,d.^C9FUL3;d@1=FP5
8=XE8N=dVOA0W7b+=CZJ+1-PP#:Y/R&;ceCS.)KWeZUDFW#9)/E7:PNHfT7QSY3X
<VSe?O+4(T>T^E3&e8&2]\<1e&<OcK/BfEMQa\4PE(beVE[5T1T]NbZH4a3Zaa:(
0=/6Q?2KX1E@3PP/I@>_PS,eI]/ZGX2@V)W3ggC1.M)@D+@+./>N=V8RGU^0:\A.
MNYVd?F4Q75bNf^&]H.^5W=I#.JdY+NT;=gadeH:;M2(YR=AgN<bPKbEBROV2/^3
YG+NaS5GTV1Vba#U2deX/<^JJO,??V.Y5[^HS0ACR)-6]?7MA#>4/=/_N&G#;;a5
g)^H++KFMMMg?L?DLQGAX=H+e=(<b^I[KZ^17T:,+PGV?/2\;B0@b8ec4cg[9VgM
Q1K3060TM6]#2R-H6;\eVEW)P76A_I,W]H(?Y(7c>\eI91=WIJR.H/FW:JU>;TK9
46XLRAF.\?(d^(>DDQY/d957:BeIa<Q?F]/NB<:E&.aT68eN-b4,Ed?b0&W-SN3]
F3<M\\++PU/F16T6AeQ.T7f2IRNQI/#0?f2.V_JBEcW9VHV94FI_R/ME+051:d4)
9#a+V9/)@T_(;1]LX0@&g]e4TbT(4]Fgc-9@RJIGAP9#F<71QFH[RC3gY8),__W5
cXQGaS.2U&6#:fUb#IUI#d_d]@D[MYY&bL4,acPS6L16OYd#I2&cOSbF5&OD:)4H
=7]J2++JJ>bD.aB?fM2E97MS;\7<Q2a?d&>&ID+P/46W\5R/JG:b.8c//9+++Ed4
88Q.+5.FKV>J1I,[^NO)7HL+A6[3=9MZ&>UPC_<R?CSFO^-Z=g1@-(48H_3(9c7Q
aB;@eR1/PV?Q>#+QD1MH^6T9;BM?Jb?\\@;NE[2&>^6I):-TUQ?/HGF:ZZ9:-CXJ
F65_^H7[XfQCg&:@^KF/MZ9=/g;R/?YLIYOIO3a^#Y-OWRU/L:UQYV>(F[?,WcJ^
VQXN3<7P[IXBV<-6.2E8U1\C1cP,A,;+JL#.P5a:2\P_>4U1e3@BU@E26+16^Y/3
:EM7Cd,U<^(47^=^=HN)HCI<5f5)cQ]M=Y(,956Y75,Z#H#;NB0,)dS\0[IdRUb4
.&/f5(0]@3Q_2]&06?DF=8f>8Z;GY_,8N)TDCVeJ--T[VVK9._B:RNF[gU0-eD46
H9USW.AMeW,+BC<ZE0Y2B=8/Fe?W@T152?5/&P8[UH>eMKBPMbeF3Za&L?_IFQ/;
KbDZbQPUCJ:bGHYLK=/:AOOEgQZf-T.-+a+:7U2-Cc;g-HOS\J-S9NcV;9DG.FP4
2L2OZJ.I[W=Ga2;d8&2Ug]dIM1^g4ZFJe)@\@@4FTdF1UDX,^Z92Bba6K^,LJ<7B
cIgXd]1WR17>Jab1QA+2Kf=^=WQ_5_;B1Q?IT]):@LG@Q,B2.JAg(OgJ<3-cE\Y.
B.d;S@A+];DY80FNC70LP-AH1/O9Q&<fP?@3C3/C&99fIeG\g8=<SJUbPW#<I<ZW
dOa:QNJ_?UK0UC3gE1LX^3Mg?fS<1G+.9^IRcQ+gQBCWCXH,ceK0M)[fP/g@,J/b
+^T(K7eIYT\9[bK/:#dQI5aPMMR(Kb,5E0<\LTGMg)Q[-<c[Ke4T+^RMV9I]Fb=M
@1B7@R72c/[]HP2+\/#TR7BT11Dc(DbaEe]D4(.YQ.JBa=WfZHM:NDE4J#9.8)2\
Sf+&=FI6eba<L5TEa;604GZ)X)XXB@+?f^NA?EK,GUb1]OYD]G?&PRD6HWSXd6-@
.70JNY1JRUOQ,#&a+#D+.MX/_:U8WJ6][BgGX,4A,V+OZJ-ca?4Ba5#_(?LA99=d
b2UL6/RDHM7Q2/QB,38LG1)ecMa-Y98074;2^LYPb;,CY=5e>_-5P#YG+24=QX90
Y8U-PX,FH\#RYC@[O(1657ePd54Ob#A9W#g^L0K3VDDPa>0D:eFMJ@,B<eTQW^/4
EG4+(NN?OY+9JQQU[;A7:?C[eb\E@B](.Y_-YXf)WT-)3W72P;Q-#?,?[Z>F#&LY
(a06g^<A0<>?,DE?.)9&3(8#5FH)B6?\+[1&?bXf<3ZeGW.J#D.bGgd^>.GI?8[T
<g5XBWZS1AL8DQAbKM.@\]FaU^M,R9=3H&EZKFN^BU=D>,N0NFXLH=,9Z-G&8J4N
4DV32/O.3AMXY+@HB<HMfUPHV_NC/=S9c8Cce0YR=0_\)f#@eGe.0F@6T1?X(KX.
=(d<ATOXPA59^c2+;OHWQMg6Y)06N/B5eAY:A/JD]KJ5B_fFPafK>OFM&OOL3>UY
@+5URG4+@[da?FC_Oc_B:c1.BOSG;^V2b53Y,d:e_NUP:T3&_Sd+FI@XKJN3X34P
AY@3+/S3>D:E@Kb5JDFe+\MMD8?1.]50R_-.O<88;N]+ZAR5X(CPL\5H5O+J]W\7
;GN=40&():WZT/Jbb@2bFE>7.A:QD?CJ(c2e+?84&+Q(bb5C,[_7[6CX>\?cadK?
T;d4W.Y\O2FP/DZS+U,EO<&G#OGfW14<#_/]^B^H[:FUG[@.RL3\3FZ&6,.gI^-d
T(7CIH(2YHBAC/RDUe@,E@9E.XB/7>U#@\f6V(6:)G2.VF4b3P.YLU<Bf]\=NcfR
U7?X/D=?UT6;EdK\V3R^1e\U>f5PYR1F8EBJJ&]8OfG.K]:4)f+MgN)<,[:e;(TF
JKU051PAGT34CPYY.e1&CS>g0I-\R_3/#;;31.C^M9>B)fS0aG<0_C-CN9Z\>(Te
VNR,daG6WTT=/SK]d&a)=2.+W>\T8)e=YWcXQ&.g4AgQT8X<L>\KPZ\Hg7#eNQ+A
3UNZ:@8F4>76,9;,73SGM5f8B9C5_20[ZOR]6.b\0L#5fb-1OCSFXe>@B->A_^1Q
MR7T=eZBK#_D1YV(W(fIP<5WDcYee8.OCG]TSMc>a>.WR-?=BE>G750L3B.O9638
;>067fQ@\V,:9&?GMO[BVZ>.I,F#\a(]OH(Y4]5V=^>0Y<\<&WF]OKMb]5)/dSV7
\N)#1D;@]XCQ/8DZNS/_B?e:M?IeFXWGB>g^](Mg-I\\-VK82EJOPg(Y90K-e_4)
7-2Z:d&1&G]eD=S4?aNX4Xad;2fL/27N7g[c/W\XBRQ+-&/MUPXP1SK4-6Ua;Ug/
@K6=[BSeC_W#MQ\]U_9HIOQAK#/=Td,8(\9&L)DZFFC3_e]FQFeG[<TDL0AYRcB;
@GR7Ae2DVT2BLN_>\A,KHB;EJfN>5+de;Wc[JZ#4LL#@(H+LF5;Ab;OD^=B.)D[,
.2DUgDZbDRaZPU8@B:Ne-[G0MH^)RcVe1\b^8]36J,cGgFP\)#3OG77F:1d--^X8
1\J&36.N_F@+WGHG?.R2EQ9[eX\;_PN7P[CG]\EBeeO,+CDAB;I211<V<WH6;UI^
G#U/5PW1<+FOC2FLA?KgTX#?fN+:];9-Nc(V9IbDcY0TAf1FYB;_ZNT=#;]]dc&<
0RB^[,AD9.FW4L/B:E\R5@@e_aaeTYDX]70bI^BKG(g)LWR>d/:ObIJ^\EDVIM<Q
(R,JE_KdUfO9NKQKE;J9\.XX6D2XGHMPL4eTS7[HcJQB<;FNT(/(&g[6_HaT-X/@
dA8?8N8F1dC;,9=Ig=^/VD/DJL[S@G8_OJL(KB.c#(X_-^L42[T.P_E.=\Eb26bf
F4#>OE5KUQF&_IE+_(1R3NJTCcW_\eW;2LF8L:ZZREHOICR^Y6F9;CFSHY:>2/(b
X?Kb_XcQ4c)LQC&e-)Tb10[8]9A_d\/^cD:7[Jef+gV]A11(L5a=aR+8/[S60eS0
aZRN5fU8?UM=Z<:+WZ??AE+c]::FU(TUE1NVKfWV:&]3RdFGJ5O[PZ#^#ffT8.C\
VVVZI3SFDW[dAS5#gf>AF&Tb608OTDQg[I+2SHc@G3(]g)@CV>B^EfM3TV/)HJ#Z
dPT10?OA/^#3_/eAMc\=:5L9H^0O4D_78-5FWT)T):@.,<ZK]S/8\_f9.AFAcW(P
,LKDEe>7V.ZX(/<0fW^HCfWBC)M,B/-7Ie@F(]+PS=IUIE23>A.<Q\_Q:PXAaDBY
[/_Db>6>6OS13QaP^8#,aZYKa=N>]a.ZG;IN>+=VSMP6_E@?:N3.]a.&@U&=,:4C
Ad8U]4&3X[;eW8)5G2ZF0g?^.4dcF-ILWeRMg3(>ZQ5=HG,R<2BL]d82JXd]>=Y1
F4DL)T?6TJc_9aI3[]H+dNYRJ7VOf9]ZDfI[aK79&A/X^OHRYEeO)NbPdL.)cJCQ
HC8g+f\+P9GS_SO]<5[1>KDa.XOYfd3&_)8=HLEe@F0(DU@(<Y;<JY(X?NO8.QbT
KU0e?4OHf#8>Kg.B)+08E;D4K(IK:-S.AQ_MP]1VaC_4\.BG=9,:-]W_4@/2(/,M
GY6.O/+;=f5QU49]-Y@[?5B)Y0JY5YH>03BY5M2:]]W8U^MYG+9He?P<;A&^81:E
&/OC/VaEB-AH]KF-BPT7E;EcB6E6-;(=D,905:01#_F@Y2d#d.5#Xf@R,]7?(=Da
C)L_IK6.928#.6H6Bfe^gT)+?)J=bd]H^)B@T6H=7[S<3>4DI&IW\]R/3<C/eP<5
eRSJNN&4.V4/VW5d(S=WIC/(,aM[fbcN<@<[4;\7JcAdE3-_J)aPI,c&1ebO/O.P
DYIW;H<+8#IX)+/=@6@A.2Bc1,E;KO0^?AVQ[8DY[a5XO&OBG3-3_ZdSEP_2?4)F
/D2dY@8,UFaL[8Q\bK,Ma#3CEG7Y<O4K0[e(W&,IWA[5TdbO>.BJIR?aU4ZF9?FL
?Cf-e5?;L@:#I/N3\]QV882M8Cf/QN\E/5UFOG?(6d\.8WT.?AZGaU]LNO.FLI7g
V,XH=;X+7V3:UNdaAW1;47cF@U(>@:g5E.;+Wg\ASF?TLD4U=P+bTF>TC6LcX+9c
_9Z_(5XZ\R90d(NH<Da0:^/T,dG]R(]X=Jbb3g[0cAC4gR-]RWa9-c;SZSWYFQ\N
b;SK.2&@;W?e][9BSKE4:M9b&.&W?NYNP+JL7/>YZ<;HHK=:c>3P(#B@\^C+e5g9
44dAO64#EPc(&:@+3F&U54ZdLW)HQZaZaBD7;AXK[T#(.[)P21a&WR#?6BWdTB.:
:DaK^D(-4I;aJS0265;^NTTD63dPGf5>OLZb)g1#:NJAMDdeed]YFGNU<>VYa>7M
I^^SY1[Y[)8E5e6GE?)+Y@<@fHfUe,V9)2+dM_R>ADHCdK0=U77aR6,)A5(5K\:O
BZ#T4HVPT63c>:WGWHU,c3g=[D2\\M<H_0F\aM=.RaD:S<SZ-WHgSA]Z5eGZ9QCT
&JVJE5S@U[P&TRKV^REBK9@^09UfAEMOTK3CHJEe]:7C7G#4@gM=Q^8Sd7WS+VR@
AD)FD+\=U_24cZ-U)=-E4>-4:.,YE8DY7(^RM;:BgRaP9>]:X]27I>8GA=/(=43?
5._UY3KcF@6aDA;5cL_LUGWA^eF=EFA6KP&.bO10d#:cW;S5V)Ob0d0(KC=5eJ)H
D8?L]P<\CGM9@]>U5/.(dMJA=0MGEOIGX45O@P9PaaHf\T>@W7V/KGG<E8H71R_\
>_?89HEP/6b&T.^;,TL4UIg,N-[H>U[ZWVAOGX1W=>5KW1BGA@a41E(^d(MR?A#^
G=(c2?g9\SP/,cJETJR7P2&>[?&0G5:(L88K><./0?T7VQO;+JJ&+XeAM>/C]MdM
TK=L\,=_U.N0OX<WWFF[[/)_I1(J#/Za]:PFUaNb>@+8RK;^VFV1^::_&A,&KS09
6T6cEC/a;ZCWcSTLA:f9XL2c.@gIQKXHT8[S]+51L:=4GI&/@COM:2gQebM,,K@.
PUX\CU(8Sg\V?gU;6M47NP<1I<_DI\eWcRB9CSZ6.5VNRGZ:_=XVGNcCe92XbAX/
0?-VR5]5POMb9R5E_,<V6eSCc#([:ZTd2-DNY.[B:9L>3QUVRHgc&;T:OU5;(<]F
@_AN7&2TfFa7PYE@NA8f#c+W5+]:@>=X>JZ5.g7]e-fMU=Ka[^e=PTZZ=Zb8d&7>
ZP=LQ[FeET<#;/]XQB9,c826Y_5Ac?f)-Tb?Z?09#CL]5-VL,=O.2=d6#:#Ra3Y,
0QK-XPSSU<_F429-5^^_XfKdeGW2V)\1RO+Lb.Y82e/>H><?T+17/6MNIG3VbGfI
8V8H=>]F0HY<)#6/[JWS(F0P)NXe]J,Yb)&</VJN]Oce<FL1:SE:Ff,\:f9WZ4^;
.=PU=#WWgQ_XQ>\@WVF6R8=4A;PNG&g6TRTU>@e:JNgBG_PJ7cLUG1L9JT4OX/[1
03@;@W/[5H_L1>D9Q:F]F_LGWQL[2aRZQ&b8/CKQGY[,+ALK@5^@8e4KM4HQcZY[
b7fFK.J-?&0YQFK1VdM8T9OEC^g;L74NfL8T\?>G\09>)--.EIX/#FZZ\SC:2?FY
/QECVZMTWCP(571+Z=b.QTB2UUU-]_6]cKP5-TV^aO81eJdZK3.=53;^dELHA.TR
9gEZQc4C>VgA=4Z[H\,UOYD[FG6EQA45W_[0[VOAB+\=V?TGV@3AO9,VXGbY<)\J
cP/HATWDS_E1cgA1N?&eL+9.)dJ3)=,/X\FGANGeV6]9[WR0P0O-:3?O#GWdZKH8
=PM9SUYNES[2O+F]&5+?ZPXg;L7RT[F^Q<F4W&I)?aAgWT\N6EOK#YC:fKe<R;+5
[Pd<>X:B>:/D/NDV5U&J]3-Kc8CZ+]5gN>cN0]H@MK\0<MZa#:]TLDO6Y@&5]^Y3
8E@g4MORgb>NCfWXY8#F84JO3I@<R#E,]/V=(K#_GLH+])Q5?XcFFdI#(Q<^>OIM
1(H+>DU_LRPKXK>dV)B@QT2?K+/61]\c)\Q+4M0gNb(,/):UeXeC,MaJ-=ZEaDXP
eKfac(Z\eI&c=NGE1Q94;_/fV(fe3aZZCOH>:eTS6NJ\ZBOSW2bcbGIK^_+BATON
3RFOA_SB:#:dTA,J\KMQTR:g7cU>G<?LSP>ST1?8REN&&Xb.@1PQEcF-gHf<_>Ke
1eP9]-f=N3U^5&BEAID-X-DC?Cb21f(T(N#79+V.\.<cFYd?N@\<>Q^e^L9g?7?a
Te\#fa9^(QG;L3P:831^cZF;f.@J4E&JE6/+L<CZbE[a/VYS<7a<8&.=5bJ:7c9T
cd,cO]1FD))M__5&8cBO8B8O-C[FgJB&PB6-OBggV,8)gVB:WIIN@L9B?O6:^@W:
Zd[TO2e8?7V/bMdcf3U+6bQO3:WWI#fb4JLg@M_DK2[<3Z@WZKAa8H9JB#O8_L<S
@SXNUPB^S;IPb58>7RTgA9/bHf11He;6@@ZQOA;a+:R#?\FS4bNQEO>a1ZeSP,S.
>4.+K@,&.JIK&SVd.<W11HGZb&;([<T4E\5bb_1GA_DUbJ]=OR(FY8^5gg+T]fT,
b#HP,GL?bZ/A-E#GX2C[_H6Q7e9:E)7O<ZSC,8@HVV[-_JX4PB)bMUE6[QQJEX)B
QU:_&QB;KeE09g&J_R^/QfB>7.-3RZXS@Q7,[EO\Q^b8V#ZNSfO+IgP:.EgGZB9H
AL2&D6<NCB,E3(K:;b#Fe08^V5(U6Ea_b:?\N21=807F50@]IR5SM]5Qa0=5\C2L
BG+4>+.Xb_Y/<cGHAc(E_(8[UUUPDbBUPU^-/M8@DS(H4B2aEfP(IL<((>?2X0)O
IaZ9NGXeF+SeeHW9B[;I;0Y??Oc_MZ,LT9HSQJZeAX-^.G9C8^CMSC.]CZ<@SW[V
0UJV]Td_Y2O_X/[F\JRb0TH:WKEOe;&5R>I8UQ<CG(NJad-<1VcbR8AFE^72A,9&
,#YV6ENM7X9K1bdL6=FMFBO\DNDJb:^E.Z\1aFCW?Eg^X2>@@U02U-3\Q=GZ6<L:
86OW_PERC=Q>J7G)?B]4_4D2&<Bd9G4g6^M-=/bY8H^G\?;304,10CRaT,JDG<1c
Wa2QCL;-7]OdcQ0PHN?0.(\+ZUAA-]O&/O@EMgOYM,/VB0,BfYH_O^fE_S+4d<4J
NU:9+\SHMd,\6g/YN>G6PE9Ac]4&+EZKHL/<G3/1fedY(PUGNJJ)bYF#VQPg-P5,
A-?fddd#6YRJ4]cJ\LD)KafGAY(,JO8ZA\g(UQb_a#FC7-J2Bf0Sab>HWHcEDF1R
#8MI5[+Sc/23-fP)V_K\_72ZML-E?4ZbZ\-]5@==(JUTAZH-C4[dR1X7)cC,3SFS
&SB7eT\XEgVKWBE5#6&>8K-(Tc.8GP/>O\H@g<gC=AXG8#V3g.Ig<FT^5:,b_B]:
bdeZXB3A#0_[Qg5?G_7KY>50Q+LHXVA-f8Y1d;eVe]Y0?\J6aG0D2(JK)a)-A+e-
JG^)?S?^a89]UPCR8fEe9IZWeK0I8,dH#(T0TM\4;/d--(BABSG+?;=bC\bY#(XJ
BHQ_=b/93((M4\XTC&6+(Q2<Rg+dM+ZM+ST]Ye3YDOg,XJTU6=9RRf_dSPJ1XQ9K
;fF@bc1;&Fg+[],_P#<56H=2JOdON-e@5^D<L^6a:5/6eD8Q:Sa43:WLc;9K796.
g>RC=C&R\)NU,A\(CJVd:+I)+FQ(Ke9Y:.Lg/D<X(9M\]NPK#HV6?3Z2MW)_ZH@@
>g?PFGM?^RI\^F[6HF/G\-99TC<B<;;,^/DVOCDQ<=9RXEa>9SaTU)I6YD]&@<cO
<1>F,,fdb+0I31G>(BWYSYaWE2V81=NDI#M)HO#3E;c;3D#>c0IS4J/^@I8_e&3a
>LA7eJJ?I@8<@6:3T^bE3dc(ZE7X8-aLTe>E:<18IKcULG8FWRY[1XF[TXT68OF:
baORBLdC8MAFR&7MPgYI\],7LId(>R3&T<6.+beB9?6]PQYdDfg#3#fc>T@M/]X4
/H3S74.6:YS4XO@-Y4McC^[<_OG]G0&2_D&]H,P2RZH9._GdH[LQZBK&B/R@GG6G
FbOR2deF8[[IS1CJVGa]a-OR1OLHb[R<03de152:X)]?N_/72KA^;)?N(LJg(&TI
7>;Y-]B.S46>Bd1I&?+#DX]8,4GR:?FAO7S5JB#FNL4C/MZfc6;T,gN+Xge2/YUV
IaCK1=#EcbM?Fcb7U;7\S^K5C(2R43L[[Hd9eGPCg-eN(TK&AN@XR;9?L1a\E]C^
dOR3Q#/NBeHP-f7Z.X@G_9;f/_HeP8WB-1eS[G4B@??7SKb&f:cWIZ\f@PEZ;[_/
(,BU_XdYeS#3\.g,=<:^R8+^QSUbZ?,]C\gaF=>1eTF;QQ>Z@(GC#?AH,EY<L?LI
E?>//5gP41,(>^71Z<g,UfKJ@5DbcY:MD11SaH<EXE6K3;87>MV<EP_&:(ab3+BH
Fg2Rf.\TV0(OVfZ6Pg#L@V,VH,e5d4H)9),+^@-98C9@JPX6V/\AELZ3OO_d>#Z;
cSPJI&K^fBEdB.a8[&]]M>#FB>)2ME3fA#U(&5K4U@@VLEfNEIHUgggf,@35K7GH
Vf0]R:S3,&[bg,TKfPJ_PO^3TXEO_4#_P40MK\@LLNYD_2),]U9_g7f]_YW\YN@G
5OV??3+NF,A:I4XHR@\eV^E<UMaGg^-/NVLS\ME<AL&&I>&+(c4e(@Q6#M#>2d7d
:e+BRJK2)96-:::K&SD3YS63@4].?7(5?,_N/C(+-gX</0>b\XGOU^\5bU#c4SIc
Ga(5R6Tc_PTSF)SUIB_MW/EP)H\X?aUOO)e\9K.M,(X6,g8)0B[,).6(d-XA(?OM
4Za8@@U31X@gIG7)<H0W6U_NZG[@O^)^D-X[/UZ/2.\b:#0G\CYaM.1<3WU^W5G/
g6B7E83<TQdfa:_U5[Z_-/a2LD>V^2#U^D04FGNH(U01&1I=,d3IDYMeCfT:2AC3
ZWF#7BM[)egZK4LK4@P6-QFW;7ba[<L_T<QDVD^>GTLU@]17W>cF_L^J<IEMQCEb
@E7DFL&@WegcC7DJ2BY5\F@TBXbL.4/#gI/=J9cKURgY6(>cF-.FU<S]=UI[5?5N
-V9J6eQ@dHg:D)OVeTT+FK>+D;)dGQ=fLD2:YDQGdCNb-2VU+0<P<1AG5(53O]^b
]L(GOSYS-:?WEDKHK\YGEf&-E\-=ZX8S&Y9;M0KW+/6@aTGg>EF,eVUbBb#c00KF
R(X&B29X^W1B^.3f&(eK:HS]T39&;g]@7VD;a:^\GRgY-,aA<ZQ<FQ_K]-/=Y,)6
NKd<]44bCAc8623>/(dJ[YDcW8gE2gZ_Hd+C=,Id_=?d-7bC>MZG,=G15a.<Re\Q
W&-;[6A9#;NB5dg=T1LY,eN,]44ACZc[X&bB(S8RPX,I)e]BE(<c.fTbE&bO2_g=
dMGf3BaKb9)d:[-?Tf;@:;9V79-?J8U=].00/[GSBJX\EJ1d8gED]?Y.O^)DIDKX
9;TZD@bV>./aQ3f4/cMa[T@_@cN#C=#<:VCX3G5F^<>\I1@2>H@^BZb\4+VZ&]:f
LO#P,_cDGCH.gJ0A8F[=-AbNbVGc^XUc3.I4^KR19+KM9F3e7cU>3cV-:SRV=c@S
H((UJUeOTL^)U8R7F)f#Y.bfJeP8IeU@&().bY4C]Mf1D3^4=BC?J)5Tgad.9g\(
J=,UAa[G-.42(/A=/STFC#D(PJ:LV+Fd[BND/e]ACO/9ADK34=AGd5B=a/)a4KC.
5E)_U3RZOJHMZ2;c4PNg0.?J,YTdf/><Z(731NR(ZFHZ-b#(UJNBQN0.g/BQ_UU2
>L&BaYe@f_d6=6]V.31-+IK4TN17>BMDf1HfL.\E/T\RT\gfNAJ;69bQGQ77D1d-
)OJE/HP/8-.4((+ZH^aPK\?X\[T/C3-]SCQ:Q4;SW.\>R+ee(d/6Rd]8,1VA)cA>
N0IgE4#cfUUB2Q&I#;aF.@?IUS]GSU/@S,Y30&Y;?2WUBY/&f)G+bF>@](8#c913
ID095Ve_@A9-FHL,MH<F:J/eV\@R\W)?K2<1#Y8.M2IgJb9@fCf)7V?0(G7/L(dD
_<VHZ?R^:?.-8247#-5GgE1D;FXV7@a/^>95,9[Cd^I+FH8A]C(f28^I[<9-B0Wb
8H(:S/D<;-+=)e0Wf1eYHQGQ,S-#6eFTVW:f3+H32VYT/^/SB28A=N3Pb#Vf]P9Q
]1fL(7,:GF=2T)Q^fM3JXXfd)_YFBGId(U@>M.bGBbX&Q?&A8VTXD_WKX][JAegG
>+:32U^<3PPKLC920-b=4E^GRN<2]d9X<7WI=43+g@?54F6:>d3@gGO8100+?X?W
WQ+H^W9G/J#&Z8Q]-US4][G_aC#CDM@[R:CSSNC=0V]NXBDRFBFB-[=GV<#4YTOD
B]#R90K/[I(0(8&eNI4X^(20IWGbg[]_QDfe0DOW:fX[fTV8gd)=f9+afP9LNbRI
e(KF/c]g?<=>D&8;VTFB.:K@_:Y)K6ceV>[.T^B9IH1=?Y5-,I\425AX<e7RLV34
PWLPNNO#8-7SGKaX:N\DKS)S8c7RQ-##6+]FgW,A7H(/\983)0]-@YN\aP]#GDD5
YC(P>#O:;[])HQ48S<ZB)V5NWeI8VL-;,&:6DUYD5X8/?O;B,]+?CaA+._I#cT7J
2TdB]K@G;<E/_(D]e9bWQ0(0Ub54<HP2f,6MIIQT4-QT>FRc.(fQB38]ZUT,aaQZ
<=TQ>.&?VVT1<K;RbR\S?FLR)_SIaaX\.GdZ0;c\fF]]&8F2,4G2-/1f5WF/LWFD
H929?C4Ng2\D,:eXS4Y@K=ABU>/YdWPW+d<f/I=,/_0(/^Y(PBg,E1e<6HSCY9(b
,/:EWWRU/_^0W9?((QSHJF,29E0RWEOZQ#aBC4CM?#JfT?.ZF0.OQ@5ZXA>FZgG=
#d@&A&aIA05@5A=,G[_2OF@;/(S,3\Sf,WN944\^0-cFBIS0CR.Fe@fd;<MZ=^R:
#1g_V7)dXP)-L,d4^eA)CD,L,\,),DbVe/J2gZ+FUAf\e&4(P_R<+U0Q_\9T47W,
aC3HO5^CPD0f^g9a=ZC4Cf?Y;-N42V.SfDb1_(]ML+&K<.aTeH54PYS<3AaNIbb7
QX=1:,W72MI&XB46=QfY3^OV.G2B2X7\A5)GNG&PaJ][Bd#.M-H]CU#UdJ^S63R_
58g.&,U>93E<2<+f-RS5R]&C=LeF@H+:JK+G6GFFCE^9;QOMHAFB?^8@?RL@(^(&
S.?dd=UAa8fIR(:@4W&,Ne#@7fYO/LLAUT(K)I7O0(McHTXW<F&IC<QP3<^QU\-(
PF/AcN]UEIXY4Gf#@8<c\?UEU=8?dIbc;,9-ed>OX.;NHdSW,H11UW7+<C@1HYb@
0SgKG]&.KUb3OL#U2@)Obd]KeIDF7=b(FH[7FPf#&4@J4C66BSaL(AS#K5_#]SD&
^O6?>XTbAO8F;IU=V064:Ng2UYD1LM&B.(?:#;LMCSU0<W<aE>W.9+TG1Pg[41]W
1TQb=K;68eKCLB=AS[O+:(8Zb.DN9O2NJ:BZE^c]]#g\;g-6BORO8<1)^YC3E5<L
(A+5C<G;1DOB@#^JLI=0=_BJEUfCJ[Fa<\YG+,G1_=cfYQ4R];E/]@O4=Kga8W80
.+\EX+(dE-D_E1#-R1<Q6I9@<0F7;bJ6Qg3(_PWN45=NBR2K@Z9-GB)4/Af^CJF/
NfQA_d1L>AH;If[5L\:[R.3D#U;gFg2A0RQP>=(Hg5@F8P?B8;(37E<&Af],NN0N
bU@ZQXMPXJcVD3I_PCdR?eB<>D3>deXAa<gD436MHB8=A_Y&LIH5^_TQXM:\^,M:
@5KF2a74gM:;4=A3@C>f5#MfKWWOd?(]49\YXF;ASI[CB8IWg^D_GZc,ISC()AJ+
CWbE.M/PS?7X2Z>X>FS\-g8d\\P3U#Z]3LIW;NX-FDQ?=g7I(dE;S@,;dN+fL2HF
T)DU??eF&F>;J>P8<O6+G/G>^+J-SY>,Sb(4QFHeDO[VP._6(.6^YU(H2EQ:CPXc
NI[QCN\M=:9;-A,H6>5G?,83)-9\#K_\]QUcgUR<0=YVFRL43?]HL:U5IL3f=5bB
89_Q7f0:;8/cHc10T32192_=d=gf_]E>g6=QeWQ5/@TTMIQAe4Xc0Za:U6<2RcH9
[VNDcUMFM10S[V+)1_F4.M+H#^DPaaR45-\#4[@6McJY(/UV6)fS<T.6R=If3bGg
_&<HL.4V?AXf[gAaXa=)Y7&RVK-U+K#eL8(V=-JO:.:>Eb2&f2QN)TN+0^(IBTP6
<4W7,\W46?5[+C8D3R(gAe</V3WM8Z9c(ffK1^9PG4+DQH@G>4B768FYO+R2T-SH
R6JIRJ8SS3_^A[>]K0c1,#/6c:E3ID_OR4)KHCa\?NE8AgIb?&B86#\/a:3>J^b=
aA+5WHMcEE,PX@\J<Q(HVB@)T:)XED3KVAMR^=4>[f^]OFeMSAMO9cM:Z5XcVUHG
6U:\U8BNUH(b@=V5,/(_RHF9\ECV]EEUBH>45HFN_S59f[L?Db2ZWdM\2:C3Y)HV
Y2W(HE;]1^7Y=VL8D#9>;;GNM1(/Wg8=PG,^>[#Ea.dZ3-U<G8>AdD/4Q@58b)]2
X&\.194=[2:Y:?Se313]ENdK+HIE;.T,#[>33],3;4SUb(f;[WP;_CH]c3YC?T+9
RP7Z_Y+I&;MIC/d=-e31+F)F?YFcARH9JeBF#8O<WK9&_8:9aRLaNG+<ge24-UdR
c^=G2T=^AF,&6U\A&#[_[Sf#1dCH#:114[:=9X6:;7KI?.cKZ>A]8JaTZg\Tc@Y?
&c&/A:e/SMaU[TI;#;Kf?>G_I?a,C:7]_Dc#,N?_dW)2L1a@/b>d6HB(Jg(-8,#@
C@)a[KS(^4EQ98J1MBXc^H<V.@+<I]Sdf76-aWSXB#d[43H/S,LHA1:\/Eg?;+3W
);^GLI,DHO:#cBPXd-P=@,+a^Z.Yg@>J5QcGE<JVZYc#aF#QG9(QYK.gK/<9PQC0
6+Bg0d@Cf//H2F#\(9G[YJO-d+Y)2W9b95M4V.S+)@H#[HgFHMB>WQ^OOeARNU9L
b<OeMB&-e8L<X/DW3V9V.@BE0JYOcET>,@WZ1(,;\-M;R?2:\>IJ:?ZTDN(]9V?H
d7J&M.a(<NR)&@d-?7F#-)R#d[#4X\5#,eF43HNd<S=W^RR?ceU43N]XK:_[@[MB
/eYE#O\2T8J\f94^U(L\O>92Z+.;_/Vc994DG\,e9&b+C;IA8J>/XJaOR[NV2=4G
BE)gATWW6MOb.79UaOD=?)B>8d,1ZcNf\G3gBU2)cQ8>@f?26FA843?e,S8X&9;2
1NN2^.=@[G,XQ<eJV\9E8OD+:NEa6/<O^?1.RHbB(,AP-ePE[.bJS6ZB+0c?Jcd5
CGJA\;[@RF==0I?c(GeJ[8I;L6d2E-Ud;gM?#fD)gd+@Cd82)g_+[,2_G=gLWJA#
D^ZP2N=K=\AB+P>bd15+6D)F8CUA^\I7>&3&,-2FWK0@U:]Rf7,8ZeF/:^ZK[cPg
GCc/<>I24)4A:dG3:e7TZ(:.14dEAK\=I[Oa==,_]M7-\HU]?9]KcdbgU=KJ#XQ#
aLTJ@bR=_gOH_C#9C\c=Y:V9R<FaJAf]0JQ0/Z0T,W.I7E[<)8U3QDD)MC=]CS],
^U0]_@4.=O76JRO(Y.:_#6Y61S9W@>A1-T=U]7CC=+]LPe6:LME,FNO&#4:PgFJ)
OAG^G?^8)GM4d3M+^-aR/gbQ8EUV5[I+(QILdV9\)YU:d>G:9>^Q--VGe&N<.]<K
7IL@P,PGHP04+ARR-OSE4/XYE#KBRTRU=-d8gE@,A,+I\Bg<,S,F7FQ[P6[&A;IE
#^Z+^&5d4_:g1HaEJ#Q[9_9[1bXRRW,&4R+-9HK#Wb^cX>8^Yd0c+PS)V],cW7,O
)QB6MS1D=@OI7X?MVNI&JbF[;MWLeY<1QK^^8BW+G\Lg\8bV=]U8Sa0bbca>f9L)
?\QB@4E;ZO70fJc&a0?a57)9PCX)Q>HKf]6e^.:]Jg/#5=3=dB_&9g\AW64Q#Q>B
UD2?=FPS^(4bVS8BaT6?&Se?NDFWD^75:XQ;6.Ve;?=?/SH)-.4,OIOTNMRM.eE+
2ASgJA3CV\KbX(@+8\7K6VdTL@FM0Y8P]f-BIdPJXM/.S./BVgaSZR=NWU_5&VJA
cZe5[be_H->KH061^\X>Q/_MdFT8aUT#IPAc=a1b5&9GL))IKE4f)<7FO_M^O4O/
\3bOTZG[DZQ+5+>R36^WF6[I@G2:^3QL(WW7ZQ22)Z08DgY,S<)+/^.^D+]dX.,8
9WFX>ITb-J=O(G8g.=@Z;E8=X_PNQ+XfOgY+G81?32\O;<(fR^M;?;e=VL_g;UZW
&=H-ZI1Zg8DV1QK+ZZFIXCcW_@Yb(+2E&D&XZAEgGfA.(IHY]0BEgJ&+1)SG<KVJ
Y3B-<TGLFAUM)?^7Wf9<a9a63._@.=cX5=@&8B&U\&-X:Lb4E,aZ.^O@QdWJH=F/
[5c2;d+J=>dEP9Z=#_8(WATLNV5I14@d?FL;HGd/K9<BSW63<3-:6]-9/NeB=b3@
@H3Igc:[-e&I?2=MX.\6Q&X4gM:J[1<VH>K_c,?b&Rd#e8f\<dbDg[/D-IX)d)=:
S#:+g1ged9]2da6+0MFCD7?1AZ<GZ3>NgL#HRE-12RC2V&8Z)=dAdLf##HURT\7=
-XRLN8KTE<[9K>+9d(;U)D,.NM?bF#O\?TNcTY:90DB#]CWO0Na@HIR44V]WFKCX
eLb[-+g.61B\?@Q52VR)OHe5,[Z[.VKSgf9?f^gf&,+[b6TKW5-e=3bCG];bLN7a
Z6Fc^SZ;]g4Ib<_(6:NNMP+GXfXRPFGH3Tc3S5aKI:X=b1J[5Z@1LWae[961OI\3
X)L&eHUBQPBR?M;4=L]+APE(?f.E@8[LXN8NN8/:[f&?XIfdP>e]b6#GI>T2I2ED
@OeENCePc-#,-[89&1E0\MO,aZdT<3FEcYdI6&4Wbe&/>7X5M#e@cLS-N5W8a:^d
KW5>DG)NA@1W6E5C&YBXQ)DcZ(;GW>H]BaJ>LV8)CgZ;YP_-:4=6cM\K6fDX=gYT
,Q7AB>D<?NB]YL75a<^9#bW=,+D(CS^\.M:HF3G2^abZ/W#H)W\CIP&bE1bQT0XI
R7&+&?J&-C:[BZg]<(cF1(9^#5JB]N9KPgN;(X_c<Z>?&B-1.=VdZQ9FgXNJ/NP,
H-HJLYSg5_SP=&G2F5B,e:-,Pa7e+Xc[Y7YD[6/RP2_T)]\gFB?>4+R#4DLF6R<@
P]7YPa=<GD<\<e,M944_EI:_ZQBTd7Kb;UWZO]@+\?N9?W<[dAS2DT<2&8bS/cG(
P7gC81[G=#0/#>Y2UMMW9&:54E?W7N^6[(AFO.N+4a(Z6/EHU1YO0E2_(Q[U3_18
<3B]&)?GMOAS+b+d9IPHDC0\UTN6KeVg+=Bg@:7B_2U;7#=B+SJ)0;gXf63>c5Y_
[T5HNM)W&E98gg;MUATZC&T7WQ+_8#-<eIaWIDXC@:E7GNS_)@gM6Ug^M+G^bc5O
980G1O)FH2Q/5/SV_JIW>ES-,8R4FbP9CGT-RU34X2=MVT:_.>3g;C1TG]OfOSR.
.H(LXC#(aA>Kd2Qc#.(R>Lc@D2ff</L.+QRIe2]07^7:H\70-f[(YE.aKS999:A3
D2UZ4CK0T=WU\&UP6E>c(98.dGQ_JaJ.aIIXSFW(Y07QF:)=S<0F)V>d[^VP;B-<
+&>5M5>#]V\OcgMPSJ4OWc,]0g<O6]E?^d<V_@S]\Z@^bQ],BeWcSPDET2VLTge\
U4M6/X(R#+0PO+c]8\ZKY#.7OU@9TA-aS3&NI)7@g[bVO_GG;M,gd\.S^;OQQd(]
3P&=KgNJIG2GgIbLP]EbO,6CU>NVR,31(5+[Da@)PT>f,L1HcNW=W\<0E?68+T:>
1-<T<D[;]WS7^B;\TWIOb_CK)0LQ:L@/49&?RQJ@cWbdg7JHK;HTg^4>TY=/8\BK
e:RI8dbD8fgDeI&dJ:<<+--1Y.^@BbC(]Cc4.B/-+XV9,^_?5RAVJ(_OMQAe/Qc^
&a\54TH:_gG5MC7_?7&a-bQM]e@eHNM;S9Rc:.\aZT.>BFX)d[g6>VK1DT.bBP>e
)cE_.a7(c:F3Bf+(.gfO<=W]U2GX^-2CcM5VS<Y^3Uf+PIN.U:6g\9IM/aU@GFKO
>Y#K^8NR50?EC8/YeX9857P+H4MBMU#?#YH(99T1Y^=F;.be8e.)a#)Ua@gb#^=f
8e991VTc[CeQ08O&X6W=B_6#bOBF)d-g+O@,&0(ce?L+<-^5d546]0^K^[JC+^0.
EU/N7+3YJ5?A7YXEP&be^UA;Q>b/89Z8?C7g_-TXP:P0-eIgU]P?F;5ZD-^Wc(8G
APefd&.U-U(M38Jbd::6Tc20/d&UUa)_Z,><A_g9[8\M>J_6cOB)OOBP6VR\C/6.
M06Ef2e60EMX3Q\OG&c::/6F,feG3P&B4T<OFXWZE?T3##YF.J38+V30\Y\3C]74
#+,b>UG[23]:K[&F+AWPNKc&:VHb>L4V+Ke6:A<Z?5QW5);SM#bCeN<LKB@7UV35
3Ke7SDI,^X#,?Fg^IG1[U>S(7]?^)Hb@3XDTb(YIJ_bZ7CLaZH#.3e.6[HDM[XN:
:_]I&ULd^6FT&.Y;WdR]VLffYS&&<CX10GFcIDDUg];c/NeI<L0SDcXJB;PCc6YU
BO]VQ<9@WZ6_7P3?1SCN8K0(IJH9AE7J>SgacW(ZHKQB>GJ+5B08C34X&LW9B2fV
94I&PF]&gO0DFHBQ9D\PM3=N:W_.0#A)_WbP0N7/X2PeL93#cQ=QCU0,C)B50;bG
21=IQ^X[2UL/M+<Q/d=J+/LNQT8O:URGb2B,+EcME-,2/[>\V0g:aK^6[>]FAc&3
G#U)W>b;G<eAM=3/\RL/W9VT60#BVeC9OYYI)^fUe6-/TbM[C[;]#9-+If]V?>LP
)Yf&dAYR);?-KU8CFNe/UO;ceZLc./Q6#:(<D1<H@7HXK[J-LU_E.>FC=+DP-CB^
0=>R)T7-g:\0X[;WZ:GYB>?4QMZ6;_7OM\4+RYb69)]?bS2Z0c&LPMEWPG.Pe2\C
3P8-g?9(7I-XcOO^6,Y&PNM4M3aF_WWOA]a+&-W\-2#M0?OPG:ZK82eJ?b^<+gJP
2PNELVX7,CIC_@cD)c7LD],?KME,4ZBgGLb^5;Z5bQa>S:W-T#0;<PSSD@3)=&73
cD[J+LbD/Z[Fe>FM7\T7XBARg2<4I]AS^^,O84;:Ac@2YG+]E4/9:O)2A>)P7^b=
4U/G.B3<I+f&H0/Q5A,&D)&DDXO(b)Q\/\aM&UYO+H3SO5:1D^fQ=ScQDaBX:W7D
d41H-R<CLF9g/<]TO.<?c=^W(VQ._JO(M7f()>X==H4PeRZ1^OENN:&?7DBN.d<#
JY)1>H1KHS,V/M15JIVZ2[_S4QgT#/g<_a:2eVNW_Aa8#3/IK?TC35fLW_M.Ca5S
+KCLY;/ZWP8U&P.-c._L7G(;_VTc/GM>?>1JFCe/3S2FKZ[-.cT?G\YM1&=2#Z\:
H:KFE<),,\G@4;DSG;_c_Mg_3W94?^E62PLPW#[E_,S4,\eec6bfG-U@6U0>+63]
H-C>J)LWJ<;gF1G9BR_0G6f[a=VdIMK0<\db_2VTC]IJK6TOP5JH0cWe)gJQ_dY4
;dW;+AN53H7@\+FD^U.7AXbY4bg@+J,X<\78]01)0<E<JRdL18f0?66N>aLZ=C[?
[70a^7BQ2)f^[O-GIgGQd5>]HG-VcI,53,[Hd(:=AG^54<DOP^>eHNbKX-8aGCA5
g#ETSQB2P<cVT1IGf(SfUFH@5bER.1PAS_C)PJ#)<W/0><PXXL0A;;dL/NKFURD:
=GK.27Kd(bPJdO6FUPE-8YScX94[J>TDD?CM/AXYT98Rd@,T8F5O\B?/SCK\B>7_
,9>RFEOU;W\F&ATdd4,W2UNY7]\ADUbGG9e),;JF^U&_9ELeNbNPASYc^eP0<7XH
[PcA9b(f/e-961B]O1A<<J7T@=S3d<5FX8FbD[gdFe01Q8<KN,YK7NJ2>]=]1I^U
T2C@EMU[+D42E2<Pd\f:?f1?8,VfQ34Abf,#RBfF4XUOZTE862Eea&UfD\/.#53]
XbbWQ3L6Se3_YeDJG/MM<a_(b-Q+-aXAM)X#T4/:HI>P]8)D[JXHFLAf6#8I332@
f_BUH]ZVJ#g&_,KEU>R,+d6F&Cd]1H.2T[76TCI:B#8XeZ9<)Z[;dXaS9dWSG/Xg
V,.QN.X(0R2:&17;#_?^,Fa5bPdDBMO]6;=dN,H3_UcOWLR\[7C5;Gb<TDZg0gH<
)?gf0KXd)RI^M;],Y2<VXaJ,#<7Q?D[gYbQ8=7T[F;,H6JSI5(W.HW(E+G:IL72,
eAXQ#Q0AN;UC7Z@ff(C/SY<J\C?JV_QM\\+U?BNLKdJ;a@=P^+6b;[92Z_J)9#NG
ROUOMM9-#e(<Ue7Y[F6+ZgLaW1Xd0AZ1dE(BMQ_@@C#.cYN1eH02[,1\X@QNa16b
&bW9cDVLY(-:gDV7.CDVH\<N.-dM<:;3],O@D,A3>(_4T#TV3I7/ggW9Q[6MQ<JH
]QG?gU\(A_L#0RdEe1H\<NSd#WH?SBbYdB<LbRddB91@#M_FU=-W:MWP+:b(^N[#
WN8_KYc&WN#=BR4)D[dKA]K229d^eW>KR+KL?=5C\.QD_-<5_cH?@<I)J7-BDZ9B
6I36?UQ>&ACKbNZZcF/SY6@3?bGeWD+fT8IK-=Y&dM(0HFEcJeW/N0J3WO4M?/9Q
^?e^]N;Ge<Hg#c]N@]?R)NH:M1A2@b\IX4(8g<=(.F,B2eB.22A8NGZTWeP&@G#E
=_:MGf#IG.;/ZSbZ@HgQdXCXH3IFNG=d:6^<2c@]TV#EIBcY6UXJ_5RT]F<FRbe,
U/(9#Q1_fRHX15WLD)IZDDUHJZ),<NJ(YV.ag-E/H,D/L7PcHOQ&JX@[.D_TZ>T&
MHO-,e[3O7JZ4a;(,Je5Q,5QbFJdA)H:gIEJKN3?3J/2da?b@;T;I.dP0bTPB8Q&
8#:K&R6>=K.M-FeH)LaK6db1O([8&R:K?.\72fgNag2C#?Ig4J@K4X.=CVZ5Dd@D
6Z#S=M#896KH@.])^5-f8Hf<c9M0MY3O8AQ)D/HeWS:0d?-25dgNf/:U0@U=YBVC
URGd=EN0KW5/+cBdS(?3TI1;Z[K-aa?IK:dFK;IE8,&ZVN1,>Bb<d)3ECfVT#Lg?
ES&c^YG5E0\QC1a=<L04fJR3P1[A74/U0SYK0-RR_JULG)-,a4eLA,XP=4\0;WOd
EHN):29QJ^L-;8c@\f<+L&L-,WO(V^8IWE-N@?O[b\cOC=:K-c<9=;f.e0395e2d
QJKZ7f_75)&_N)L(;<U6XE&[^QO6[&E<SK36UA2G=.0J.^Nd^(gO<1g(OATP1dOY
8dbT?^?^OaQ&R0G(_#V][UNg<,4<cXSd\(LZ3PJTL0X^,4:FOLe)BBFG:cL6]cF(
C],?9G_1,eDKRRV:Ic^,WX[_FTIDdWSWGIFgeKWXbaSUFL-B;);T@TKgC;-;afOc
PCYGf2g<]b[S\C9H#RKXP6V5]bD2F3@E:a&)g<#CgF[VPD-\JKZ&/XHT6gUg=0]D
JQ1WQ4<:Cg>.ELH]T&120?G<]OLg5OFKKP\M><H3><d93BEec69@FMeEC_HOAQT.
]LM0+Pa6[:EM&A2[b:8PJbT>9Ua5FfV55C-/1Aa#R96-Pa/WN&&+RUQ0TL-?G=.-
Z/K63N#FZ8I&VF,5\a+EMHC.MS.QE8(V38Cb_c[1(I4Z;4A4A1c,WcJ8e-F)Q[PJ
HQHD4:.NS<B?7GagX[>AXUACVPGe_Uf7S#;@L9X;KeY296:D>U<]V4S<Y?5Baa&@
UWLVSFE=6&;G4XTURU<Y7<4Ofe_Hb1FFUS<_?8M)_#3>aKHW<+5>HU:b[O>MJ<O=
4gG=)+dP.KVeD^DF6Hf6.Na]GNRW>K@P^S7]:A@H>P>f[HJ14OHPZDQ7_MdGNRBI
U7=6E4f8P6-.;1;>;P]=(AILDLbYT?1&]J3;MAZMGe3-UWKFI\#?g6bFNg]9GHLU
,O2&J5J#EGHBO,[XFF-0+YFcTB&gQ7-gW)H)._,^g[>)bH,##,MBFfY[5MD;De^9
fQM/OP1WeX74Y&G8[YaJG,4-3I^5:Pc6&>g](J_(0YML74>L6_3?<g4Y(:ecHeW>
RV<T,+4GUE28;ZNOL&RB1=&:4G&(CC4C+8-DF.\@/f1RJ@beF&&SD:7RgL[?_YV(
VA0WUOXAVT2MUQEF^^5HV9P&9^#D^Jd;Q5PMQE6&fW_PD.=\D@:N7GP/\T/IdG&(
U6_gMK&K#aD[3NCN\baAQOZ/OS:)QH;L=eTEIY@;9Z5S[WK_,Zd[/@F3AGeTbVS7
FAH]Vdf@G=22-<X41XU8[S)f]VNeP&[Y8(_1Q,TW[<eVG:/\#<TT^,OX@(S6:2TS
A_2_Q0:^bQ0355[X:JN0/TD3,3\0gQTfW?T__T+T^HE)Me:QH75eB/[EA&#7=1Db
2Z<g2J69GT@A4O/IQ@-A]EBHFJBe>>J;KW&=&R8CP3f,K+2a2/M^0U_^)^\\;9.&
/P?5#HY9J(Z)3Z71H>I,<YCNdFaJ]YQ>Q5-9SU<_Ga\OA@:)DgB4eKSaSE<aE+JH
f&X#6R[<Ke9cCQM?f6JN9c_+B-WA+<V&49g,VL/BR[b/<e-F+ATBVY(EQ\>BRVSa
ea8?AQKAOP&f[4M&][g.[JRBBdX7GC/OH-6.Qd/BJ-X3QQP?E/R/TNeaUX-:&3&A
,HE?).?M@86f5C/<<?^Cb@GOJf>+bW]bgMLB<93cJL3:MAO]IFQX.NB6I>9Pa66S
;Qb]A86YVTg25H+PU<LE/U&84QT9O#bRV4PBT8:VADg(GQX1K34-ZL)#F^ae2#9g
,B-3O_>?[SgfgR,@@.IfANK:S#g#C[/=\]F6V7=OFc8;-Ib-@32(\3@I)b_FH)M;
&AH(YWXGK/>eaF=POAV3LDg=7P/.&)g0c9J_9O(6ecYN&dCQ8-QAZX9b+PdM:D=/
#3FY;3F[-:M]5V:^>QNEKScJ^0M2D=5JaabcA1=^B6^(O?6P:8Y#:#XMPL1;S/+8
#\f09;;bI&H^;1YEc?94UW4e3cXV??B5FM,27FT]H-2EBgVPfNV8,(R>6Y-Z(dbe
Cd)_c)]A-1Ff:(ZW<U,d)AV9gP]SK@-P-e[V#>5S9QY[<?X&FAO2,.HQ#NOFC#Z>
RF:I\ZQ\aTRW6a2;S(YJdW?>O])UAf3P0Hc.II3ZXcXFY^]d[eP_A_[UM^YQ9(e.
F=N,&OR4N)#11c0J8-TgM&9AO6,DAJ+H),;(I63Se&Z:\S[-1OX/EfdD:B)04e:U
gJC_U[LeG_Ba+TK^P]aC,5=bKA(NQG+C\^3Y89-=L-66d75\9WZ+O<D].,UdDW>\
S7[Y0>KU/DX5(?0T,:GRPL90T3I&]2S6:B>&@fD8HZ9NC=>JO1V5/Me+AD9T<?UK
[;d0c<\V57Cf42#I#8#N(5/3_gRQc^<Rb/SG-WTR1[6[X.QR2Xf9DBZR4)RS-8D\
GdO1fIX25+F@5\I7VdP:E;c^dTGe6O;:^aOI]@K6@/?/C.R\+a/.de>;@VZQ5<D[
b@<Q@J8;8N^7;+(D+\YJ^=B&-e.CcR<:aL\=[@64<&O_,YS^ER07f#G;67]E?=>N
-0=1#Zf0Z/.5@<I0Rg.7.gXA(_9O.6d2M:LaQD0dJV[E1(aERYE8.HcOKUI(G:g=
C@@0009<(?JfQ&e_3f+6aLe#6)9)aT?HfVeHO^0PE2B=;g;7ZSPQ2=DcJITD6KJZ
&&7e50,7/QMB&3K][(?9KV)?1^NH/(BKQ754VWX)?3cL)X/0/9K1A5<^TMdgNZQ4
Y5>_7dO;/CGBQ7[.eK_cO@#NJ:,57?ZF.,D(B&W98#D.C,bRcgMQ_OMS-cKg<<6@
;]#;J4-[-6T\@H<2Deb<MggRE_DT58GZ=M#@SSX)[J\NK<\X?Q(<(HX^ZTV#F6\V
.ZcDeSVA@^5V@7a<\GIU7d26-P^94AW_#>E<+.(R;97eES#5LCM&:QR[a:MEA^@2
TEL-_;P2O0NVJ(A1=F(N&ded^6edR,d4+;NF8GA7N&TG3)bI4ZLb(BdJ-)/UR<&e
-[.?8SQ2CA5Tg3fND8bP;#Wb9J9KbW^9L]/Jc?:7==74@3Q/Y(cBYRF].\f=GUA7
<F;>;UKK-OO_L/D:HK00NP^]PP0AR2J64?dM(5G862@QH)S[J._R@LZ.-J2OA;_H
3<NbT>V[P@NdbDdTc<CF97J)>;M8WH46BI>I\R3^6D0>4^Wb6.fZ9f8NeA@RY26C
?8g#.e+C.ddDc>6_Sa)YEb.LXg;gLZQ.U/O:.b7d>SZ))7g8N.PE_^YS\Z8gd#&.
3-9U34#?_3>2FGdC@3-(63g+H1Tc.,b\MMUEI2>3+^RGcF1.Z,RJ3P?]0155I.]b
C&89N7eM9:J8M\JK06_:U9g58=N]C6MF(Ne#;M3&B+N?dR?cV=]0J3ZY?/HS[TLa
e;Z?8XWYeP_^geY>U&#U,e#8L:Z,Ta?IDa)d[-QD-U.H9:Ld1#fGQdYH;PDMG^G7
G;ORL^2DN@[=ZU=(5R#ddXdWJN\433>.5ZcPWCf[Rg^YTAPg>^H+dH/PW4P1)V)f
gE2YR4H6;2g,I\caZ4e>IVb5OIXHBCG[?5c51U(ATQKQFG71R3d\VX=WWYRBH\V2
ABYP)&2NL0B-ALHVBHg3#,K#Q-6eM;2+MX<OA<cOIZ1=geYJ>5HDMW]c,be6MEO+
.b=[c<7BTg=QYTS<gd@?gSYa&4KP24-@,cN+._??X)S+R,8.g(/QHMeD0cM?3dLf
<1e>DI8g0Xa&7EFAG8>(8C^]D=W8TM[daX8?bX<@Vg5[/:#6NSXc\R2KQd;L<LC?
0ZMdI4P6g/6+D5SV8L.F;>5W3,Q()J16Fd,AaWO#d=-E<].0PSd>8L4eYEPEDa,G
Z9<>76?cf-^+)P[>G/P6>^P4K_L)+XU#\8b.756#E\b/MQ^NP;ZX&1RFAN^&B&aN
_N5[XK:;T3JGe;Mf(d2?)D;^(5>1Q?,dcC7(^P6R)3GOeX=gC\Gg)a3ea+M.:fLB
1VN&HBfNCIHLYY?.;JW[WB61Z-+_)P?E6L7#AWN>@a-S<B^gO>W0^8BZ0Vd#eRdX
4,acT/(F,OC)7?GTD-KCJX@EeaI>c6H/&MHRDU;_(XABQ)aWZ9,:<g<T1VJZV<Z8
=[\_(K[bP0CULN>c.KM;Nc>S-[d;D^GgL=:UbY[[#5AR5G?ICb:fX^.VH7.307[c
UEJb4c_#WD]-,).F>g0OW>A_5N7IA=7+:B8@)dI:e3L>6ZUJ;S=XU3?6>]VF:,ec
N+PW@,2Xb,S<CS-Z?QR1)>@;J-D.8NI[@D.-cS;/L]P0;&?^>D.B_7B2NWH>;Ad)
P0;&=S;XRB_U-bcG1ZP^4LTS(e>g>R6d/F[L@INXGNRAeX7?HI#:7[fN&/BYH_6C
I9/(ZfYZE]B5QMP<g+/X]]A/=^T/#F]ZV@eO&151,B<+L9CRPR>;A.P]_X4[+JOR
N^]_38S]KJSAZCJbTJA:PG_@5)ZD)dXV?T3>\c;JUFIaRF(JT\Ub8.^9:(JU1JN;
fXNOb[X;-WZ#_CY39-E,Z2P2NBJ;L3\4MgQA,bcD^;=Nb@e:X2:4c:7P52;UeFP=
?K?,dQLW[ZYZ7_N=NLE(,CBM.F3HZa_8@eg1,-Cc#V3?)1f22f(:1OWJKHE,9b::
]SK]YI2a6a#=:<]+EB-e3^QV#Yg_,@G9S(]&+>:Sgdf0b8c,8c/7&3Q=/D6,c8+A
aF1dVQJdSWA1E:)STQg1B4F2HOO.\)@/T;-\)SE<XA(KILBUU(Re?T#:3Q6E1L4:
L0\W19e)U2:16?T8>;M9FKW:>a73@KTa[\HbH3#EPK9ZYPI88d3cD];^P;[XcDK/
&JJ-VK8CO(RJX<DEA)F>K6SQP7N3Y7;3(?QCYF1_V]V);R2\d55\@d@EH=6F>[7]
8gSLBe,1Of@S^T27^Q,ZZ?2+(&5L32/fV[2HNCO.dC9/9bZN(.>S2JKYR7&5d6cN
;]P,[>^97ZUO24ZF]/VB/aRIJ.a+dd1=&,:3YV=/+S\;WQg5a46f45W7/F(2d6EY
eeY5)2<@]agL9gN\DPbOK]DHH3HeY>dP-4VTP+1:,dN/b2MM\a1de^f_VNUf+3J\
;f_bFfD+cf^8EX=&:)E70M&.EfM5W,QZ;.)4Y?@[C_Ie.c>HEOYg>LP:XO,YIF1g
I[&,;]ZfJO9,S,W&[_cJd]Q<5.g.+Q1_0)bZZ-X)aX55C8bMZZEYPF:=4[-KS2Fd
e[fF.DM.HZK/YAgJ-MLgYM.XR/g6^5HY4:G<4fTS-&J=[]WL]+B9=AAB[_<R&1VO
fCOS-B55g8UaW#Z3@YOSVJLWH+^+^I?_82GKH7A<1P1c[Tf@=OG:eYVWWT.73Q2R
Y()=RG(J9f5KOc5N[Qc<T:KXe6[KRPbc)@DC4/RC#a_SN_;F2GgD0(9:R@B;b9,<
#EJAEV@TW>c4L:+M6],J;<XL:6]R_eVTXTBMObR08NHeQ[e=&3SIHd\=Uf?15KaK
bK;AJN;DVYa5S_[0J]VK\W;)d)+V>g[JI&)Wd]>PY@@:=SCc74X[))NWAP3,LT:>
LAS2TCBJ_##C\K_fTeBBFP0,eO1D5<^N#[X?[a(;.A[<<5,@2W^+(eT&-8S5gK]O
0b-62ITId&[M-8(V@Q95\(+7AF#RAaFC/G]@6L,.+bBB1@)JE/[K/;e0U;^45)+9
#X@H(bVHFI/A@YR<Q9CQ^#=/fTgUS9/fE))4XFCgVXFF;)Z/=b(VeB6EL<X5;DGc
JV1:RgK<O7C,@B&[9Xc,CYgC&c9fOM<agW+<I4c1QP;.)X.\Xeb[HCMSFYW-Z7P[
INADO1X+DS@7,8N=5@#0;J6cX(_Ke08-_.-b[4&1=ILCGdbLMK=@&1Q-fE6Id6c\
UMA].]e)V<D9f&de4A3=)DD_[g+R8O43.>;B>9/GDIg9^?.,V20,Kc>P.,VgBG[D
IJe]98(<X&8D^f29GCH7aUf-+G#5?0(6PT?,D4DL+cFD1#M[-Yd-R\fK.d/aQU1J
^HNKYE7N1,/S&(</T;f_2XWe+A5+#Q4:@>gA=LE:[AU9G0EQ@W^-^++(7,B>EW#B
PE5B.L2be94-YHM:]39\OOM=NIIgd_5TeB&VNgEE@3^/7AEV5:Q^P37g[PWLVReN
N9I=H1HGE]=\FT6-)Q9+01QRYKe:@bXA7YG&+FDU0]LI8CcY[7#/<91LJ:5J\.]<
^7WI(=1[_?\bOJg4@JV,:U9>,MdbGW>MR2([c5V#9G;BV]aX]A732_OE/;)UA1Sb
5[WMDR+/-.WNK?;@4.LZR5ZF]^+RR>;QO0]S)ZFWA-:<&4HcE/dPE5&c@&FD[[J@
^PX3LW]VJ9=3EV2^-4^28MHb6_FC,,BRgM=3c5AAJ,D9E=NC@5@+8&gb0-X[95[B
NZ99]]3<M@UKRg:UF=J(]BQH;LRLYA8cPOI&.T-]M,5:2ONX3Uf^cVBB-YT.dNEO
#P2aFRBOfbI6X0\RZ\]HebG^J28gC4E[/FH8fL67W2^^\>IX/7-:GDc.Q1QV#6<W
_aNULOI&Q@Z;)D:V5M99GEGGD^F5_S_2AU@SgC#>42Y@W)RVI^]BcNH_AHH.;Y9\
#_XRHP_fZ#\3C:O8S]_WG<PHDK-=8\4G+MA8+MCJbTTS(,&K66cW+CbA68]PUB6X
(U\bTE?U10WdRBRG2H(8fB:;G^+U^cJ_0==VK_J;##OYFRAZQ0)^OAH#6AQQL5R+
A3M\3NL2=eZ#MJ3SB9gY^?WOd:SY7^?(TaCUd,WA72_,d^JK.\7E-7K&OB.WVU_b
@JR,K[Ld&MRU->ce_1&7.E=g4HTNKaVF91GF58bQU\1aGZ_(V<D,N0#bXg;eC4bf
F,/8J#Ee6=@YL-?;QWQ91>,-db<ZDO7-VCJLENKEa6FaY:74(XcIE,[5(=(Q(?0E
fP.A]FNUKdXa9GUH(C&#0>]7.Oc[gLC2#0g#)Ze77L2cd7;Dg/?c[2@_,LX<]5P8
HMF_2g>U>22O_c,I9aN3A-O=:TeW_aZ?)=0bZ^N.b+](>+DB[gALG0WVa;WI.YPW
a4>RDIaX>QF/gJPCGUe,;<-F.H507_H&Q_35B[@aX8X@R)<4[(+>ZX&&c18RYSB7
,B1N.<DgX_XQfOF-1VDL,T5Q+g.[N1?GQYXTbRc+L5,ac5JX<<WHS]C(>\/7_/PX
@,,1)/a&?MJ_QU=-fWE,?K[&O-/[+U_2I82K+&^E;>D_/I=?;47eb^QA(J<ecW4<
7_HRT,#VBBfLQJ4Tb5Mg><^6TRX[FRb)5?B9cM?N,=F[CH:B/6gS?9[\QTgDVN];
4Xed)/g0,=f1/@5R.6)5<Q/AVHA1#5^3?9\+:GH^;9H._:bDU?W+f;IOgX+?0cJI
>_Y0R6H7+#ON-g&N41G_OeaHb7H/^772N81+aeLXc38QfKNT3UO(d<M0-[BBRMNY
W0ZPWKVCX/OW8Y_Y5aJcRPV^3(<,<0(6bFM+1#271MA]?BbPCPRZKIB1Q6YJ+>5I
;Va1\;34]?C(:ZUc:f]9_a(R#E>62)e1YQUb;KJ(89a&RGgGP[fd)cB[X7(G6&Lf
\?1V?0A0(501_SFQOFBQ+d+@>7<>[,V-Q8SF6)NR]N0V(c@:_X;A^K-R]gVQ+QGQ
]IEY4P1cH(Q)?1G3ZdECEX7eX5O<.#W<[\AK4VF&/,[5[7E(Q/d+L2EYaQdbJC(&
Q>f3^9Q(d(R:TOZf11DN6Fc52.PETGWXNa;a=XC,&KR6RX?GSc;NO[5_LJM/EV;=
]#,F5SRFWY:Xdd0^,eI3,^9gDNKQgF&L>^Xb52f)L&aSSPQ)a,E]fC.3/Z0@A.Ze
8IWU#UK.\1J8<Y6BN\<PR6&aXcZ/9)McG-@(fRZUWR3dUEIVTX[dYN7bdVJE98Pa
E@@d/a2F/@+(IP@KX2/NSUF<KNc0MUX)b>KM:]U+<B>&SgaSJ.FLOI?aCH0,DY9F
?F]FJeGM?A]DJXCeI5E8AbdZ:NX9BO8D86P2]JWYAU@(9^MS8L3^AV;^BY>Aa,Zd
\VM]d;gV;#adLUf<&7.6,;/6gX60RT+[/X>[BOTCRAKGK4/2]6\cKTJ3^M?#D4a\
@3G2G/E^,IJC=[BQbbe=Hf./cJgDK9B?TDT=ab;c&Of9A>ISUS4WN/KV<CGb[MB;
W];Tg>V-FC(0>588+G[<ER]4J9#ZC1C:_A&^^>3dLgJE4TYER#a0UcW7)#Lg3V/2
,T+)=\>7U--e;.-d)\d1TFee?+a,^:TN8<T0dKGXJK)7L@/;_aZEU5@(W<;,07W[
+9AXd[9@L+TM0+W09&O+-Z1]BK_GaIf0FY,&[QC4EOXDb&S5<<]^?5@:1Q+<T-]L
;cVD90X52\TKW6g^<@<E#(,#8R8G9UK2Y5#I4C^W(L[GWbg5_Ug;ZF2^80fI+\35
<S66K:\7(OUPfAX97O<gEf@3^V)MO9X?:4>Lg.8N(0X9I;-YZ,.VGEY&C[;J(=)X
:9#/N)QFX[P61dH&HT8/B+#6@8f^Tf?A:GHd@U8W3T;RWK.M6JSBR@JEP]VHC-b)
UHC7>cK;I=;O&<D(5W1+FI;?7#+N=1&VcB56A5&@[QdIV66\6:9I]a9DDU[&6>,4
a^&LEM:.<ZO[7R3D#\T./8_J:VG+5I4NTOJZKDb_V62SW8U:WUO.PNIK&aLe<L4[
\Z=UaILMN5P08YUd>DE?PI/43C23S5\baL5[UZ_S\0a_QZTf>I?fO\&AQ)VUR4Fd
1gU-UCQ_,33gMa)DYS&HNU:fWM>TMd:ZF4bZRFG[>+FST/-:5#T6?JOC71=&aLVB
:T/BNgc9K3YG]^G^aFJ1.3W9d3.e.ACR-Z</8B;gL\,LIYZd9)TTA_EK7;T,3e,.
^Yd;?.W8>[B_I6;CbRF.V_QJ6\I3@#;7@gBe^JY>M9LC[VZY)B26XNbECe&Cd+D=
C_O>?Va<F;aSNc;GMe,22Kg/R2O.gCTV/&C_=JOJ_\F2C\9X;N5Y>/I:,gTH/[=b
W;\OPW(g4E0^(bUMcXFY0BK#XSeY1ZT_>/T#PJN^:4>=4/d(=T)&DU3f>5-@\(1&
0++C@K[VdGW+7^(LbXf(I1d-^CY9f_.Sa#7G4?ZQGUB]MD-VL@XNaX1=5>B^=V7>
OUdOJ@MYC&PCEf^GZF#]0AWY30#&&?X51-E^7BeC//M0DAF^,b4.#CMJ(I0W)OEU
5-IMaZ0@K<23@H,E(XGAeg[Oaf^4:Z&T:/<+9H\RD8/@TQ@8IKD^\)OCe2JHBAb?
S8_1ARcB=\-WX,aSH2IgVg:>)0(d\9K<P:#7?7>(fd/PV6bG2#-]&#Z0@/8GE=5B
2Y=Ge>GQYeI_ACTK3_54L.0MXdZ2:eFca_d1=7@;+2fcT/GUKX=QGWdCPaC0Y-+A
:.MXL;34NfL-ZbSUEOA7e_0.[;=//)4Z\a.,;2S_IHH+1HcNSV(;c9()W&cM:a39
J@--&CdJEbE8X0YUKDDI&U,3Xg1g?GYCKT>IA,M8b)_)gGf,4;/b1TP[],9,a0;Z
EJ:#2A7gG(^HS2_TFYJf)WAH:>#,OcD#Bf(RYY#1MAf7Ce<Ba.NLfMDC5@8V\/(>
fO(]\E;3B+eC-W(=7?c.HC3&7;PJV7CK&##S]gMP>CMG17d6U,_/VW^8]eeI+a:N
U[XV;IgEV^8[WZJJ)>@<[ZE@\?D2M]/#2L5A[:dFH>gS\744STS9=5YaZDU(6=R.
)UJ4CFN[J9a5+c^=9(^J&EAGeTXI?/fWgdZI=.I.OIEU5e=K9+BZH5W.LUA=aH?]
YLQ>=D(/Z-BZ+I[1T/TBNSc@Z]VSXNGO[#Q,&^+_R[?1QYY_g5F-1-,8HNM&7B,A
Y[2\LCeLY02G\L&_F@FB>.Z9,UWIKS[E#3geV3>a@:A)\3N\Y59B)>4A(LJ8[bb/
[-Wg)?M[M(9/aT@C]aFV+A;CSTM#ET,H6B)#E2OKLI(JgGRX9.4M;J4^3d,T+S_b
ebLgM144NO_a@9ZTe9Y4L(5D;8-+HG+(/Af:EeFO#EBPA[>4D_]@6-)SKLB]^X:J
F6D^c&)7_)K:Y,;=84BfYdfNfZ8LdBOYJIE=,67EP^Nd)7aIgc9K7W;_dWAN0BXX
Z7.&_WOF(Z@&dBVaNV?K8+Q,[BeeM^PVIe620/Y4a<3SAV[Db^]WMed#FGV/cN,]
^HT>Q4W=7QS\>5(E/[DSJ70J#Y>^J=1G1b&#,9DJ<d<T)K@bY>R4I#:I[YA.H63d
RGaVHZ^XD41KX<4ZR55>PJe>4<b?R4]O,\/H7OQb^-Q@ddFbOH-O3gf(M;0FPEAY
VL,PcKD757(^EVc+XWR>7@DMKD/b=S&T(Qa^N+^1YCZ<O]F^@M9BI&A,A-YDbWFJ
(@f<K_0fTT;L;DM3KD85Z@N+#5[:,@JS3aUfIAV:Z7g/1DE2FEBDHcW+VJI\\<#@
]60QIFQ77A&G2EIa5\84./BAN=2=4f>Uf>Ff(B2_GT>]\SA.5>2VV06<+>R[(IYI
+T<9@:M.2GPVNS9BBA07L[A6:7&;=D-X:Jf>D;.^[XLZJJW0WE:^-=7#BUFTB6AU
ZJb6aMJCHMYF@TfY6_WN2.6\Y.,f=6;R40<_T_Id7/#?8RN29YX6;<cQ97CG[6=]
&Q[b1KO/8&?5DUWTBFcZ9=g=GXEG40-GM+KWRTZ,Qg:AQU@\COcOC\=+X7PFRVZU
VS^1e)S]G\/87LF4B(7/:L,7>IKPRO/9,e>W4/b[DdgYZL>I7460=;bWXOWOM-.)
dO-Nc-Y>?M#.\\@@MM1K<[)4-Q;#<[B+,&BVYKf,e-@bU7;.[;63b>2<MC24AFF1
fQ4\-7H#FZG8+Zd]+3COE0P/5(ZgLA(@8B5BdQ6cc[#UM-WK33V\^2&BF)e-2VAU
d1U-?;1A2:T6,ONEBeV_EUde8>V=+XDbg.ReG84Da.JLO<MV3W6MR3Y7dK-H)+O?
^HgFH155dXU;=B84:V_]H>+b&@F5:;09#=OC<].GJTY3M7G]4^/f(3(K-^7@_T0B
-2,K@A#PMPGH8L.6,L=OAR<T#A87X>:G@_JY)JFX5T6:G[0,<)cI;^;(HHPR4Q8X
e2LRK-KcaSbK:&<9=-AS3/^4?8I-ZD</AcR37G8D>cDMX3C<JUAZV_ZNQ++Na9Q2
79(BE9_;WK\ZE[48<AXgD/OQI&<E9ZA1JY#L5Fd0eMY?+16E4[a?@2[RAFWTR\]2
4_<]J.^:>5X[SgZFZbO^GC141,G&GFIB+H3,2BN<:2/PI8TEPa@2fBKQ>0/=/R>8
a;Z9g]?YC0WP3&+-eL0#c4@@9HUg(ZY/R2Rg3Q0c#>3JPW37+5?M#NfEO)92;eSV
A^C>TNg=(ZaLF&8/TW-)Qed,##Y-MOJP8fT43X]-B/g.FF\/FbK@^ASa&bEGBa=G
]CD\B1aQJT;#3=2]TVWa=EXWHA20KI(FG>(>A_>YA)_CI9MY2fUQ9=+f-K<&VBOA
[7,VLY5OdK:&ZFLDP=,b)&;O?-3\&W[S=1P2;49]=<)1&&f0N1cV4?:&e(,[W:12
A@5OXV#5ZX>+L<eWAfX>^;LQe[+<8G)#CE(g_WHgAER1N7T@bX[TINU/D<:(ZBL2
4&_+1=Y8LQ;,c>#+be#AEA@&E,P<KPfB,Wg_5P[-/WME?TH8Od@:N>6KMU5)aES+
5561WG-Z=Z8&3F(b9GM:>?N-[(a7=,IH>FOPJQ1UB1d,75O.fM9[U66\7-bG(T1W
>Rcc3.]2KH5gC&FY)2Gb]_@gB\9>CY)YXa#/5OJ_@YZ8P<U=:0]0^X1g/&@?d#5X
\>5KB^[#.fER<I\c2fdE26;=^(#SMa-HZDO@H;B.Wg4<7L\SN9RSLSd4+46a>H7Z
AN4Ibf4[5CU;D6@-HBD1F_M5BY+Dd2=^S;\6B+I4.&+FPg/W^C9<.BI@EX<Y\NV5
,TF<>Yc&BD[64-0?V\H\1OT;H.>H800dW94#@6g75:[62VB=O_b=>>\fb#.^C64a
8IcME,XN@NSaaZ?ARa5O,>9C_K[?a:(TG/&gO,A#G_e[T7aaMO1BC:<XD]VH=Ab)
\a=?6g>aaKJ#(LB/EF?C#\b)NUe1e,PGaWA2HL&695;U(\@XXD1)0VI/E#Ua03HL
J+?3V92O7@^V5c-MCFST?>P-e.LA-Ta8]86&KG,O?Fg1(BN_9293ADHP;HU7GeM\
65DA<@\UKYE/PO+#[b&V\C,+EZOI2Ad)#0T2:/-gZ;a5Fa/]8JGGM<5:,YO#W:1O
KMO=HM)0dg;=5(ZfC#ST]W_D2?aGd4ffAK0V.Nd1I1FOL=OHX#MPa@)bMfYSHXIR
+CLRRf:V&DTf>,5:?P6)YG_C.(1a[6;?.OO3I04/E8N<dOPNaQN:M530dbNF.^#B
4c,6V>WEA==I^QFe7O)2]M6c[N/0W)4g7=&dHHgK1Q@f8KAPGT:Z#UMDbF--&N1)
09MfBE&OV/MZZT1cX:9]OCO4U36S>V,=Y=+LdJ)?ZI1a#+HK1CZbC:]LR-,FBUG:
?T->g+AeG\0^<0F.)a5D:X2[F>D:4,3G24IRM9I\5dFFVPS\)@Q=X<b]L#2LQ7-/
QJ2b?T.8fg/fF#-8:]0#HABcI^JJ):TGb2Jdd8aeI9fX1QH16FBbFD>YDfA.4LaR
#J@\b_cM/7>G)BCQU[W9W-R-YAg8\S.PA.NaL6_M>3MbHGCKba=cVGASb^[H=6f3
^..?N7_L#Q[IH8N37a(4WD-d6(BeY8Hd#K_KSWH#M5YXCQZQ?UBH?)1(9gfCaVOf
ZU4QHYB(MF6_;TbMBAJNQ\/ecc3L/4;aSE[a)QG;>_HCbKe)MTK&;J6fNTO(I\A4
)S95TM7^/ZFD:(UI=[2Ue7bPM.8T>;1RK7g(XgaIb3IS>,AD<M5:8K31_S9T=6d]
c&0FA3d]RM?db_W-X-T=_23KFWY5\COg/8:;F0HC-eMSE+<)TEIfB)PMFgG]Bd&P
S6.,If0H,OZO5V)CY:;P;7MQ/baM9+b]-_X6:9^beE(_V.]#./Y]/e8VCQ5]OU-W
\/7N4I+)6c4-AGNWeK2&OIILQaKfJI07(O/,.P)Z[KO[]WFPV.=<[]Keag;GN8;Y
2gW/VO+HIH=aF0^+=/gC8J;d9I]P<8A6@#4)8B7NCC\7TRTAFPJ,]_a:6(O:dIAK
4g_JX3R>D)2E3[)@:/JA0aZ2<[TIY@OL:g?FQ+/#O&A><1>DZW/J_(>0V]J]_;5<
_</[K0E8V-4bGVT8-NFD?E+&?TJ02D]fc_b+a9ZgEd_M3T>MP,<M(,\Za6;5(0;)
9@Hc:F#0IUTXBg?W]\9NJOGb@BXR;Z3,41R6Faf5F,V[F&Ka#DVbg-6YgZL6M&>E
F4HK[JDJ\;G^6?X&dDL8b/.dO/3=S1[DV#TEI1]F;NeCJVg>]T._U)5CE1]9>\SN
0W=>c@_LL[C&8T7@5]JP<@J]/6N4;B&HeZ5V-/D3I(?N#Z@/#+,6<37:J9RZZ=/d
e=XEF3VFHP]]RbGA0-KQa].BDg)CM6Ea+_5.S.UV6K[bGY>aJU-fd;Ia]+Pc&5OS
HF<X-NGH;f62RS#26]UY+9KH5Z;LT:.3fGS>_cS)Y?^0Ve2(WJ?)BH):=7T+)[9F
1Y,Y8?8R2I0E#a@H&6SYYMP0ELZ553NB-Q1=-]:9\MIb&<BH+ec?6UABaWT2e/<J
PE6S96<-[ZVHW,>T49[UdY>8)L]H_-06_dZPY;WVV3]C=:/N5J^MU/4c3QE#NU/0
-;cLBCbgO0+d7^=UBVVLdH9-INOg;c;,?b5_JI^1.gX_I<QAe--87dA9F\7Yf2,/
\(<f0W3\P9/>KKD2[&MEd,LOe3;bT/cbH22.faeB7e(XNX6CDNR6R1KX6(&_K2-R
0KWN(^1P2Gf2eb=W,Z(:f03b.D8-\0bGQ=&]S,J^#Lb][0PZ9fa6AU##&DGB9X61
7dg^3b/_COX<Q<@g.<&gbD@&5WdY66ZT-+PI/^15Xca]4SbR<SYa[8++C)I9NJg-
10[Nc)>]-[8A^G/;OS:GNH1d^@gJP;_XZ:J8RHGVM.QQ2G]9?W(S9-F^73GP_b1N
c(X8_))YL6\eZf=fQ>Q4=W>2(37GX#9[>1G47,<,OU8:7=b-V:?U+GeOTKaGfeGF
L]@XBNQ?We<?YFbPddf>(9=Z7W-8TYL4Id.4E0cX(SdaHf&a?[C0VU;4E2A5a^7X
P9(Y3V@2b@(^.gP#W#>[ObIEF3?#-WgRY\:U3^I#/RdED^fZFZ4;PHb(J>N1TV^e
+dDWKN=UfIfY+90aQgKN+?D@=<Q(4=C,C_)E_.Pgd<eO@[[\d&]9[)@OaaFLUEf<
V?9MBgLOcT;MD7X&=S61g)eZ7PL?SO)7G_A<c+_NCdH_^cOaD>?CY,9DW:@-Z1fD
Fd_[,?6UX_^@+RRdZSWH]XRE&#BZJ@NGdd-F2:X4.Pe#4Cea2(M^?g>J8V=X9MBZ
CcR8e30fgd,^.Aa]SO=\#9A5bFJBH.f:f0)VA\L=B/d0]7R,E<cf<JKT>73S#RII
H>J4//ZL1-gcH[C.S3aQV]1\SX+Gd8PM(;82gF24+fUL@^#C0O33,<BB3J)U8ZUC
V:>d;)CK[TVO+[XbHFFWdBJ3UR+]#a;J6[=LWU\].)U,fc.UE-N?_>&:,AB^7#O\
;HgK8/DIO-1\#_5](eg5CPFZYO/c8D#S;8CO+H\9PF:1;KDVS/&/(PFJDe=/G:cD
a7KB+<AQbT)>9b>/ZKJ.UZ<^=+DT&IJA0QaX9NG;H]L,)a078?C6cUeb\/.eII;;
M)b[23(OG37@g4N8;A:Pa_.XK=VC&0@;@ZY&J:WSgG<JH7RIf:_MZ0[MBO72(dVV
:Y2S68<IZ,IZ];,.9#97I),E#4ZTM2&Y0YSD^R17U/dg[M>@G-=65f.NKSB,ZJ:J
D1EgC2+&-L0BLG2HYNA;e,L?VJ3FEJ,.GPYD8>]]4FScWXbLGD7_/R[fFY&d/VdS
Z##^,Z_b.agNM]J(;E._\).45WT0(0Z05W(JT<<:#dK6R0;N[X&B5/4a[])@CYaM
69;H@?L417d]OdE[g7.7L:S1565)X<UfV/77]PJ>F1@.1^XS8V6)e22D1\=_OT/@
Qc@P:?-f4.<<I^Fc0IIT\4K>9aNf4#5]#Fb.d8Xd-C;]4G/6#cP/UeLY,:W(.-CK
c,PRO\9B26U)F_f/;^6gE:A[#2-?J,J0IE<;>0)[]-.2Yg?.QSd\6=f#7J3.3;K<
U&[\QKfZRe=a[aO,3]If@9ACNG>.4?GU6QD@51b/QZF#RI@(]:R/Q:]1N^ZcNCCf
0M3gE(?Y6L]F-.f7Y2C=,XT4BA?e2Y_P/_E,=U[8O1F&3+@HLAF>UZGAgQ_1TEGV
A[+?3f2OV8?HQ4e32-:;M/?N^b5-X)D3Y]3^TAZ317)SAOfA>(\b\H78<LFBXaaC
@,V+6>(TVA4&Lf370ZY2IB]7R6/H0FF@&CWQFF+dG3WSGKFLON?/()WPN/D7CUFE
T2ZfGJ(Y+X7U:PgM0I:,[:Y-W4eNePKAKBXE5W5a;&2V?]N:I0T](>2edeOc?LWJ
P9Aba4K5X/YLgBg&?JJ:741cCHKD:-/K7XE6NK6W&#?Z+LS/)8L^9?cW\G6^Kf+X
M,.&42U2VA@L?a/Z@Z3Me?a)MB^/UM0<Kd4-@]J&1/W#V:fIbU(E(<,=GZB,E]+X
dP@@,/EbO(SQ9(YPDTY;2]C,cYZ1?N[XI9#?RZGe8PGNEP,\M=RKW,F)XJ.A88>>
]21CRCKT5T&DPf+,IeE:eLMfKVZ>#AT6=KU9?X4g1<f[ca8^0I_7_+O?0)KOO_41
\H8-FZS5A@GBRd8LX&fQ>D+,]9I9)VOgN.b,]SBgW;Z@D4V[B\-Q52a=AC1B@\M0
R2,NQN#WZSZ3Q/Q2B=5D0P<=..773cQTd5=ZK7gB736aNLUR1+HJa<4YL.L7L+Ba
PGbH<.]WHB@_.<fPDM0F4]W04(QO/SW]Q(#b3P_VcAc8L\52H2VeVB.57@7c\N:c
2bD;ea8V1&dfYU:2T&^0Ob.G9?IB7gR,MV[C?JLeLbLU,1,J27P?>?=6/XRTGUVB
]Sc98c.,c)bfe5H,?RYOV@,deM70NDaFed65MgM6fL5<R\3&6G21.Y5CS:)g0eO\
V#QeY=\YB\7-5+NXOMS)AWXP\/M&bVcQT<_+<4:DW8YQR&XN:>RNZW^MUB=3e[aQ
fY?A9+8d.[,7Re-FKCQ(1.E+TU;4#LBf;KfKTO7SZOCa49Q8XNS/eCA27GB?1b08
H>1P1Y-EKDg+1H?.EdO]^O9:L+Y\c&a[e]8ZPS@c;f>=A;6.1X;6M#b-YM);1;.g
BK5#gC9_U3)/b/EE>\@J;ORcKP+(6/eX3a+f8)UMAU3>)X,W8R8EZ]CSR>Zb?R1?
UCIf[/]-fe>SI3X66-<g(?QN3:/a;gc1^aS)\eKFY=N;B:\;[-=AHVO2A(6Pc4GC
1a>P?+S(7WI=C1_5MOKH2=@P9[1N?K,=X^aFDKBMX6bH_S]@7adR.M/[YdTL_?X]
(+_G\3+&B0E),55,bAO8O@;5XK,BOe]</Pg_aa3CJ56B=[:0cU9F<L@X;;5J8VA[
R(d#J/]>WAfWHBE6=eUE1MQR7Z,JELc&=B,>RSLH_(9W(deP,.8<#8f1_V/A_VYP
&.GdNc81/>_d/;O?V+,_U-f)IEDf7UD4N0H?M7,>EGfVSf(:f9C>V=MS>Y00:RTU
1\G9\[67Lf4ecZ+TQ^/]bJMJKdN?6F>e2IO_/^)ZId:DSX@J8B3(C#5^0^[I,I_d
@2^<T_)ZIe1afAX,@R8U?e]J==P[U99FR:f+fJ&[ZO9_<?5b^F2T<R\V2W6-4\eZ
;Q[2+GT)I^Y4L^K5EdQ6GT?#1[4Me+GGI2ACYdKLYKf8E#]D?QBDGDMfRJ^aPeN(
caQDWK@:<M0B:LC1[_]f0;a@>#FdF9gc3(Cd80EC#GV_YRaS@IQb9ZdO(Z\0^W6^
e0,,IG@Qe>I^BW1a-954bHWDUT8\J&DJeb/+\VZ5([I9HURC>>;edC@O37+L53^.
_WP=X=#6P@2H+fQ<\T>Z,URNPBECP6^e,JUU_#/]N,)^d7\+a4>:V<+eX:MS/T@P
J,)B[SAPH&E#N^Cc?DX,c(]\N4f?Q/OYV@&7cI9dKdG1?P)R,1ZfXW\/f6gH/+J&
8Z+SDeFQ>a/]-3^9U<BegZLA2T0QD)>/_9(C4:6X?Vg+FPe11&(\H(H7ab(<YAb3
,Z6^&0--B0MfQQX??0+JRA;:2c,-a=K0Ue:@-=MfI,VLB^5:NG=^TA+CPAI]0Y&:
AJ5dWaRA_Bf10/QVb5X#EU;b=7L,0GaFg@^a=HT]A77#9T1YACQS2-c^6L94Z5S,
]@gbZd.F?).9?&g2]R^g:LeO=c1#KC:B8JNV>dJ?d.]-&5NDLfRILU(@9UC)?N4_
HM_9=Q=N(SKU@aF1\f#a)&P(BL36TBN\]2/aYYO>2;\V51Y5(9Of]B@RJO_:BOXA
K,1\I.5UNa@\OKN./X,;CaROcd73/dIVZ;1YdK2GB><:?XCU<M)g@U7IcC>dQ+J=
OO0E3S](DPR&8],_Fa62SG_D]C0P)[CA,S-YS-<Z.33Z4-T>5S-&:/EIcY9:II:1
+eAHTS;dK2.5HXAVV.R,K1F6eVC)bgR993gRJJK-X&84?U01_Vc_Ufe;\G#R.MgX
4\?b39/)/:g77c7C;PFLNBV&LQI#^BVMT&BFZQTY>)(K&eC4bRZ73?+E39NKc4L2
J_#:PB(7,O8@@N..1]Lf-&G?ST14&6I)7HCdN^dfBE?TO./N\BS\E:Y)N(#),>/S
3,f&0:W2O@E-O.W?K4L_K9Pc.:EeF+),d7e;4R)(\TcO;(7;+R-K]<KNI4>[KQ\B
WUb5NgDR)fb#NWObb;W@)gZbX:_4_b06^ZN8Ea7+.Gbb/\;9aT/agQ)J8eSL:5+<
A;A6\:T#1CXb82FG1><3S9E9WddAMCbE9IIC_O)cP?@Ze,0ZR9;)&A2D/1eK=D:b
7ZBC-@Ned3G59#NRPb.V7[_6G#_]396+BI+2P&SUb;.-Pb56NA(+8@cWbeRXM<@R
AGI2D3Z?\BN7+LR)AOO^>9P0\TSS-5G0WHaD;<TS_6J901bbTW-&1SR8M7:bLA:.
CD1>#U]4L1FcU]1PNbRPTH>NIbQ(^NN,J^TOTS^UJ_SgfgSJ3b<B(?fTeLDL(,_O
[Ff_>Q[]B\(O;AH1G#7Q_G5-L7[M0U4:^T47,EW4IBQP^MZce-:58U,8[EOI38B>
VY0,_d.G3:3CM+:If,S>IM3OMaI:;A,4VO0ONG2.DYH?a8M60NDg0C<:8]DWEFS-
g_7+O\D+?+(a\OUQO-DC;BA7T]4XIG#MVd5Og7@5H&&RI;CS\BcW_.U+EWB7Z^=\
8bV8@e71,;2g^2I4WU.<&NVTB3Pb.#3cI<&^DNaT[PfR74f_X0L5][DUBV@+/\Id
Ef7(.G(Z-KaNGYQP21cIf:Z+Xe\S53F/^YJ788?9<GLQP#A<[Uc;N,OTU^G/f1KA
=dNB4:]]XZ&Ab+P2AaT(^g91>)b5JXM99BDA&O,>b_&,O[?(\g:/HM@:9G4?P1.)
&).6J^Z(GDFXQL\aD,IQXF\<b+Q\1V=0B-f/?/(g/YTS_b>caTEW0CO#K@T?B88_
[e+17R>2Ta<F8/B7E2?[UEIOb42K:Zg@JBEM4;9GT;E>#;QP)<:Te=\QQ6T<?TCM
EV(L3?#=7-#f[Q>;H;M<#O=BLW#HB7&BJgYYH@=_/-SY>=NHQUR<)YaK\(&KBD5Q
#c,RZ5FV>DVS@1aNHPe^BN^=UFCL;Qd-:M7MDI+,T:JVS(OW;UGLD;CU2X&[L80R
G:EEe[,;^O]-+7HdPM_Z,Y-I,BBdOeSYf6g=#>_F]]ReC5WOSS-fW<EUR_,GIXVH
>]6(_M=Pd2d)+8[a?=[^<\<D[U_0)9@_]5#\G??RV8M(4TF\<1EQ^?5./;P-&Kc0
)R,2efM@_d-M?3UW1)e^_EV2]2[6cgDB1XK)E;>?7HOJV7&Q/?\bF+=6ReC1+HQQ
LPN.Y6&;6_CZgF(cc4d:d6WQ4J,Y.e+X<1Fg>SZO9SU/K&NB,]/BS(<TO.8(&eDN
a,X7:4g>HF+2/c\aDA_T=f<O7?GQ_&B<G&I695Nf-CNNBS,g/V^@,6E:=/+M\Y1<
/?T4f+/5_F1XE3O,g=P.b6,Ke,2R.@2#=)LYJ##>RC;/8>6/gdJd(c@L\;e8AQ1U
[_:?U/aKPVETW7D0_7aMD(K&F(0=@EEG7+Y4>+6#7E&eAV.-U)STY,N-U)TY/ES=
SfTaV)A4>QaHUf2ec0FK)BIC_\BD>\R#_3)3,;/D7IIZB9+02>>Cc-8L#7H^N=cC
GT#C)<HIMXU(;gI5N,c44)\LPH3Z==gP=2IWJBgdP>cf]IF_SI0C8(b<OBbR^#F\
Ff3KXQ<\+Z4ZM^/gSA+4\C@&(+:#\&XgYbR#0+0)^Xd7Y^EQCS,W?9F7=/(B0KJd
G\LZC^O(8gdX/J6P8Z<Z;dRBdJ)OIE-6UO43HM2Q(Q1\ffBOFIgVY=)Q5Jf)[+Q^
CQO#:MI&/:#7Q8\T.d7FN^1B]6#]6[G1YU0-d8b0;XV[fYW#O@RV+/gSVA//SPJ6
E>3d/b^=8=.4.@BQZMXD->fO?a2YYKf&0O:GUg(cHIL\HK=M8\PfCM/P?SAO+Z,I
ZIZ9bARaL?1<_TRRVAUVcV(F&9J:H@,3YDQOd_GV4X\)6aIT)X^/MM:Ba>TFd>J_
=H@S(R-:fbL=8DQYF7>bMSf&6&Ab3?\eb+OZJdD=?E5I]Z.DNcDG07>HAfJR41+b
R6H]H0.6A#GAXV;FafTLDX4IFDeOW>P(?0aK@59F8WZ>+\6d0\L#4Y6<1a6H3<GY
aOGUOLD5\8KA]O]D5(.F<c/OV>@gNP&P>2US+@>I@\F)[FG08acMG)Id2.KKR@AD
c5f1BD93\@P_aSG]e@7)I:M6-KIAJ./PQL_,8DX293NBALLfd8H]ELCXddgUNT&7
.TFKF)PB1,\>6(=)ZL?N,K_d7I4SaKfbMc3Ed^3BWG3b4-P_64],?D/3g@0E2AY9
X-CfS2]#[5cVGB@W_[7CCg:6Y\UgD6_e@&Ke:F5a0Ba;X,J6=P[T+N.:/g,+U><N
.^#dTQg13M\:RBW?T->^4c\SYHQeZ[T3V>U.@2,2]b3;9IJ[b&>_9I?;_]C@]ML(
32YR6_2E6;R1G9CbRF+3c\MY:7OF.fS_daN]A>f]0VGHDUggWX27C?VLa=5S#82f
,1aH_TOEZ71)Q@gCOEFM^;UVC#11(B[C\J,:Zf64JAO\P<5UgOgGY5d<d@B7TS2@
FGDQBJ<=],>eYLV[TBK\/FF#H&@D.S>f8+?fV;5A3YbHNB4DYD#f3GJQG(E4YC(Z
2YVE-Z^c+S(E4J)D>]5S<UOQIQ)-=-=CC(/=5XSM@SP;23f)g/SgG,QKGW+N^).,
2TYeKS7T5eRZ,+[<^8G[JO7:L\52H5T;FS-:3aOc00H_Z\LQ_8NNIM=]2:+gMDZS
89<:;<]6&2UJZO-b]]@-3QB\32J_fTM8ABZLg+Q+.4&A=(\W@E2G-(.a_K9N3[S[
\IPZZTV#Na1&Ja^5QGfP.,1]T#.K]R?bGJ>MND3Z)]B,);Z3AKH61E@_AW^CUMTU
H\95c4^\A9?-QKUH#CTIEFJ/NPY1_,Dc,0dOe^AH1/=/UKK>5+<Q;6c,/]=FaX/:
CQIXB2:U#V+WEcHIN,b8./V;?0a3WSS.VD#FY:cT=\?2)1EYAA>QNeL119T/K,?G
eHDLD6V13SALI<<fU)\=c(<[>Q/Yg(ZIfUDOHH0U25=47/ZS)&?<PVW(P,^C-X+]
_FBaG_Da7g+9L.9:F.59F0Q<TS9D4gR7HQ=d9?#@Nd12;JFFH?AV#&R=L?;TR9<c
G09Q1)eFK\_5E=WZ&ZDZ83=AJTY#fO>JR:f6g4WVS).cZWdRc@-d67&X]bWJZ(NI
RJa2@_6UTXT?3P8ZZ546HL9I2/DLCcQaJ:VYE<?fCQTc>C@_Pc_Bf+ERP4d:[e-g
7]AJg0[^Q9]<XLOD.T1Q_ZMJWK=GR=E:F]d&_PKd(?cL;?fM05.GG/:^3<72(c=b
T-cR12E.;6:&?0#_N#BUS=QNO<ecBQC4cI:F3B#7eHMcZPX[W0]N.F8ObB-9M4(:
FO@^;<]DLP5]D:H8TXTa1Kf^2D&:EXK?/MS.VWD4)d06.MEU^W[]J<ACZG.fS7PC
B^@K;Z9If4[gJ.0,bE4IC2YG&_f&dZVM8TQ\GNIBb>S]Z,3M(1[W5<eC+Y5O.,Eb
;S;//.\LNVK(+NXd#?PE#O2Y<T=Bd(:9Y3VE3E_88gFVH@(XCB?:E/,=B(B9T6/&
EVXa;?=AaTSRd/fV[T/J_(Wga]Q52-#T(_O3:d2MHg[#KHdA&S_O+:,8W@QXS;CU
NF]Tc)aAdLA=Se#_:#8E9;d#3g]&8XWH=O;)+GZ(gW/=f](F=aT:A[R;J#6QI+_@
RNI;29bZMQX7XI\dd1:?2]d\eC[=Cg2^JU@K3M,]dSP@=Z2>[+[_bZ2d:gT#b;Nf
P8.>WT)gZKBB#/0FJ3NcVO6WAJ808b_@aT3)ObcJR&U9\B1?OgH8C1X,Xe[]PN7[
>6Y=LfS,B9Xdd0XFcfNVM#18(M+=f)(54^@Ke_+_-URYSWefZTeCg6M65])MRY4P
2K/?<8bEDRa+D,+B9LUNeccFH5(R[,CH2J(LJ<0(X:<5F\L1/,ND=3L9(D^_#C.K
Vb-dL&Q]7#b(+ITU8,fSKXMM-WaNOU06J-=#:7aJCL.#]]JZb3OgS-_&Z?<^.SFC
BIU<2dI+_)=5IQ(P+RD;#@cd93=X:W3DHZZ=0/)303bOc^4HAX(dH>e]6^H#NN-M
AM7==08<+(-#bU?cD7K4f)BbYHXX)b1>ELH:?M\S+:/#-GI=M)W[ggXARO(AfcD[
.+M/\;LQB,\6DWG@.NR-+3:f_,<@b9C2Kg7QEdTMeP0gKUJ>JE7[AZ4b^(QS?Z:=
C@PHe/AbUF-14WNGPUc@U?ADB9e@\g1O>^VDD<=dgPWY3+dV)SG?1\E@Rf?):N_0
]W3gQD?^)3_e,WbJf#V01<ZS<4:EV2eK]Q_2,0Z_JP?g#O93S3&2KccP3;GL/Z#3
SS>X;_871?d;dbE,+6(X&H/cJJ4]148f4R^:2fXP\/;S)73\?+N=U,WafH(?,OZf
MT6eXK5R3egDX#b;,_/g59Od)V35YBb@76,<fN-QfC>]I6;U956KI:(@G>[dC]]C
9c@,&JD_KL+8=;V.b1<C(AEP[)F2+ABP<D_<c=Y8I1:.Kgf]dH4[K1E)NPNZP[>\
.I,.[K9eMDZEV,;/@^TY@PA,S08DEL&d;45^+/<#^&3T]FJ5X#8I7E,Gc=59\Q/8
4bUJK=Q)_KG)4Q_QE.Xb-WOP3>1+4&=1JFV)RDR3e#N<:P<MN;L6a3G]/KgCa4<Q
[g;[cf)aI?&W)]@RFH10+E-DC8;APR-KC<;_@fY-32JE^^@TP&/]7cDG0Z5a85)/
SKZW-D2&4VUTgP\_Q&]4\8S=6]H5B[\9P_WE;WGVS?-Y:BLA)?Ha=/X,9G\.fM:U
8X58]XMY[2/K^9N)[cXD]U?KC0]3:_S6Ac(5TST:^CfWa(Kg04f&MD0La4&7d2^1
?7]L/\>-BAeW+]18eB+ETRCGE]a,NB;ZGR/BA7OKX@IAS\J78\QJT_-^KB).4#GM
_N(.Z&YTD]V@,4^YSI^U4K^-S:5H:(_@IE:_e9DL1WYQ<CZf2D3_[Fb\ee>bROBO
0:?5ZL+(#^c(Z>.7J5&.H+VKULBNIH7ReVbO<>II0:V6^BOf&a.d]WJdML3AOZa.
O_\&<T/D:eGK-3U1#AfEZ]#[_XZ7Nc0U,#.0I(P/R-c:S.)UDJPV]BC)eJUY:Q^?
2_#IX5)HSfK5;I,[3baX+D-K7RbY;?+MbGN2T@=ATH)5MgVK0+MD\Y?I8Y:<Md_B
Q(+cU:0[BNRP_^agBS[HN.M^B>)g(C?1>YA\LdN&,eHF,Y[Y^ceFDK#e8KPCC2#/
H<=W?SXPEQ@8,IHeTb6f]&Z/+D)MfJ&egNBZb1)K]ZfaK7#BO31dI2[.?Z8R?dL3
fN)UCE-SEZe9e2Z_\S@TH3(f;Q\=OO/&]Z;=c-)f@E8\:KUR,(ZcP12GAQ34&Tfa
LSc3-G5&]_-W&8abEJ,Ca67H1c?W1/LaFLg<ELE,\g99[#P<;:a6(Y5b<V^fQ8W\
3RJ0@L2b8?@+9@3GR]SI3@f3TMYKM_gPSK^U2b]A8Ja\3-CF<Y)#3Q[SVY;C?JO4
WA.\6RZbESHH8#0Y>RTKUH=P^W,,J)4G<EKTd_M+.W-@SY6b+)3_Me2.g/gS<Fg,
43B0(9X=16DZ[;:5,6=:[bB_#P2I]_PbZZaN^V7QFDI4U)\-B([FeE<<@?193a)c
bJ=T<1Rf7.3LK_da^A47]Y^e:F\@VY.?fCTQ)9O1&_2#-1ZPIGW9P8[];I-@-DUW
CG-.O\30(1=##A4a(FFHG/;JA5(OKNI_Ng@6(HUGf4JG3cQ2VOHHLRL]WE+[>:Kf
8?]dU<F:a0^YZbMD@L0^/#9QPe-VcRI(;O4T:F<B:gGM77IPVcEY]W3PV&a[MG_)
JHJP]OHM_X=a^2D_^f./90_25NcI6(51Vbee&gKe0XK5dKAKITdF;_Iab&AH\YK<
\C2@ZV^H5F.69;7/YP?,HEDcc1e5PfM1@1?bQ3OY2P9(dX3YY1+V-ZR?01.USF0f
7.9[P#HD-DLRac;\-_7#Ff&@;.bRK[PI^N#&8dfd@Y]HS?IJA-e]-4/F/8YL9=T)
b5T)EZa;HM<[ICN9=[5H4_@2[#899=Ad7&Ed[SJ8T^Pb5f&NSD;NaL(>DVPRYC<U
M6EDPBCGe0D^d]/fP=Z+ea<X-fD>4LKe62W@GI0+;)dZKWNYIf4d5CZ8<),Sf/W9
VE@/[HQagU5OK347/U;SH[+2f_B)V]<>.2LD=\^5)=O9F#\YW,f3)3QS]>#XG(?:
]O-3A+YB.cd5<:<V38LH-PVXdF:ADOEA7ZbOg8?.[3W>S+XgVfD1:G9U\4MC4V9>
Q:9@JD+_4aJQ]UR(S#SbC8-XJ1Ob@(R)#fR\__>_Md8/:8N5c#JY^V/C:#X1[gQ#
LG<,\T7];eY>I\6D/OH=&TXeg.b/C>CH67\A/\gaM@\QPW@I]OYMCF=b+Ma]R?Hc
_5g8PODDRX7_SL4QJRQ-9TEW,;dCA7_<_g]A=Ba074\[d[CHL16KDaKBdC.a8AHE
H8?RR6=Cfg9K>WX).ZB(KUdQIe3,+].#[.7VOK\:,WgYY6;8+J)A#<]@297[A8I.
a16f&_BA6G0@P.X(SR+2+JKb-7eDZ;]N_6#__NH^U1<<HEgRd:4SJT1;b=6X2]U@
>K#(;_=Q@2(bQUU?XCP=O#FFX+f[a6)]_ePee27\71&SZSdf0F/J/FKQW[E:Z-//
HND_/+L/MCdCV8dQCbS;<BXA5GKA\b-187,+=)([CP]2Y@A;1D;WV19-Y?6a:U6#
O)8Z07ZcFN3EK++#7-VB1_,NNV,E2;Rb<?-WE]S.@S\2-&2ZTL[I4;>MAH=cYaGB
DTc@^f]/QFVMH+Qffc]9^S2_8FbgJM6;\8Y1]>5D^7F0G2b5@..F@1=>>S6O\\[L
_cKP[\,bHRZBJUAS>SL0USaP+>)AT,F\YHf=RF6]M8.B2CD&8cHfKKV59[QPF67H
1MX=4LWW,57=MKW#22S01Oe;#815[;8X-eBO,G5GP_ZS;NNcaZd06Y4UAaGX_<;?
U(UG>2;@#&V.I+V1J&U?\A:,BF0?+0Z[=N[@XXB/g35\Z#DAEN3fA<-9)7+d/Q8c
;&9L..<1BYYG8QL-A:)e:[OEAb_[^^.TI9#J\E9WVX<ed8L?N<P5A#7462QWNdDT
VY-a7OZ;.C+@&F2JC2\:fY[JIP#--f,O>CA2J:P>[#:H,+6]Ef,d3Y],9e;:DN69
[4S<88Tb>(F0d;]\d-&0e-(gaDV>(CA=>];bKNW0@5]bJ\Yg&P-Q+]1XW6f5f;TF
5E7#cRe7_F#;c&2AF.Q>G6Y8D#>M3T;>5[5>K870_@d9TN3\KV2-Y25.-5a32F;F
?H0,3KYb#\NdDZ7SR)A:-LbJW]H^(0CXfYcXBGNT=RI7232fYFC?,&ZN^2\c&fKX
N9:P8EQS[WI-_M7\R\9IN?>6I;.RRA1L;M\cZIP2K6[g)?3/&6URUSZPI^T&RcgT
Y<?N.H7MLRHdIM(<:4NfL@&GD,9[#-d8g-^c3WK8J=6WW@(,bB:+Z<e6>13OO(>F
W^Q6TXY&2g4d(HHZ+6afdE_bZ_;.S+[,fO/8PC.I59(?9_FU&GJ[]\2Y<A-D-4S,
cOR]GL;)9gP?04JLc>,Vg8=I3[3GPVW[_5;IL;Q=.&3:ZdRDZ7dSgLT05]UDC=KQ
7^IHZMeD1.+/L7Qe[gd^(6RQ9-K;8E(+0W>ee.D54^8^I]Z7;e<T_Zb<gR4K_8;N
^f5^4bTCU8V&N]MWLG5-M0K+<T?T[LaG@S0^65#=g7I.X)&HCG9[LTJ:LeF<AN-U
5760b@g@1QE?/)cA1g1#DPH(g&0I)ed6,#bYDDAAPg\cG;6L=72+e9P5@3A8LM70
5ICNMK&^>WGM8ND5+C<Y997XcEZ8UB(4_8QQ#<VX^cW(1])VJ47A.G,UV42Y-\RV
LTRa&KaTQ1Y3\Y5I7eLO=T9bKd8L;:;:\H?>KY:ANWT?SE1c9)#(T.a5#SI:Bbb@
TWID>..0<1>=f;=HDYKN_PQBc3=6FU+8+[VE1Oa:E^+OH/4S=0B4BQ-\[Y\4-7fH
2Q.64TA3c1B>C]3QIUE/DGSF?940&)<5+8F3[7CW6@C8d(E41G1SJ+g1Q)S,.f8B
_c=&694,C]\B[FfKI8WAd2-=9YdR](CR5XF4\BPHR[-d;G/7A.g:gDQ^7<>I5[+X
MBDaZ:=b>8T1314MAO>egYFJ0S31@7>WH\,=@WM#^SS:1R?9R.@TWAgZRB^e/W^W
F:Z3Fe=N=QZPb,TaZLK9d_79)@U[B9Re6?IH]HOC]X0AO^3Q]4+L,I3BI<_UWD4Q
>TX^#aacG]W>M1Rg84AU@MI[.E?:T_AUL=^@LC8e9]<4(@gQc.-GKE83VMH@0BE(
]EWWbG82UM+YJ2#=#-R+S,CG9a6T3JSe,[=N(fbDQDLJ5f)ZO?BZ#^dEEJ8U8=.T
-[bNP;3_eY;d#]_3OSB_:7BWQ6GMH1,Z&&VBd:_=;gd[/ZN6O8Y1/T.C\4,?g20I
8@2+8>eS+/BaQMbJEf0,X.>Id9Q;Fb>S5[M>V<I=FJU<Df>-TS2P-CG)]I&3T2b3
SY2[7RG12K,2;5-a@1.=P#+VfPZDNN]?>PHT3dUAQC(\3c[5JO7)80Da6_KAIIQa
OBN-.ce^\dI2[+V/6>Q,&T5b,RK=)7+WLJJR3G0H23/,>UgO,TBL1-]7ND?eC7UU
/8FHQ)(MQ0#@&ZVKOb]CZMO;3S;:]JSR]EO,-B\PS.HVWH<:c5aSZFc#OZG@X6Vc
6<1C1c?3d/H<_D^M_NABdI,=Tc[_P1903V3;K1:/<BE#R/Pe:N,:Q+UaX)TZE<N(
Q.V==W;=bP#[_f)4^&C?0Y=U?G;g2cfL(8f+511=Ef3@RL2@X>HL\Z#a-4#,GUFJ
Xg#Y):+LS@&>W\O2C@aD8:c?HJJD,6=>M[NNC^ONBC::9g_L;M]c1+1560N[ANHP
1DH&_X&g]Z8W8+Z:I_FW;TPG]U,KFX3UDJM;CW,AOYbL3ObB@RTf@FJ/a_1[]^LA
a=^Mb#3)gJLYZE=[5=#T-J?4f)/d8UgFQ6C1^4T3^D;f=_0a6+J;P4\;P]b?dcXR
+?Vb4TEBX=a:YdTV_WQ_?&+UdY;R/T-ZOd]0P@U@;.H_/NGVL\a:O>46P/R^F8FF
bFDW:M<[)GHRN5db;4;?>;=M@)BEW-E2?OZW?](&O54=f\&+J[2cb^;Q)Q0M?.OX
<:O<;?&b-P]C4>0#-7<88HJGB;V?CK5FeIS>PA#(f-<UC<96XC(0PR(@NO-Y7Z&I
c\b1gc(36a=BaM+<]9.7K(MAR6];YS4@D]@._?35e;8?UK+_UV&(Zb5>;N^EK7DT
3WYCTgIL)>\@a:_G(U,JR@4MG_XBCQR,ZXNMO2-XQAbAESJKY\_RdA8NJF-:DX8=
+F&#7GRA;N#MX^QSaB#?[L4&9B.Y2^W,^B<?:Xea0+\UcWN@M-<E80;]>JKeG>=2
^[O+/SIQ[35De?-XA/eZ6W]4b-5<S7BQU[LU+g.8S3,IY:.O)_MREKAWJ2;6,IbO
^(P+N65ZFW2L/Uf>_#&L^?IQQZD:)1RTSH?P,Qa/g\J@#CCYddE_M&-Kf200)[&U
,>D\YR#6fM0g.TN_]R4OG]Cf9H0YQY9=;[YWc2Me3-&YT</.0D3.a[H8V=],&@ZB
>)VaO#H(#L\Uf6E,3QO43/\XLc9V=,.@P8,(P\0/,L@b=Hb#FaFR)9]Y-_J9>&Ba
M>(/=AAgMZ?@4,ESc;V)/R^]8(e@VC]c_C\[[B;)=V@L06QXH)>C(5bc)4bZ+3FW
#:=SPKL]3:+488U:f\Xcc=aR1T=<^Q99R7_OD@VKXY1b2Sc=:aW@X>8K-VGM&fAc
KW__2;Se4>64=)024.V5IY=K.0S,\JOJae#,YT4CAZUAd0Z7#.C0#8ENI.=R1OUD
-TR^/PY@@PMVUJ^6HbIG;c<Qb0=O&0_Xdag#_e<Z>FAJU+SYf4;7)T6&6/E&TX.R
TYJK9cZSf/J:4N6De[JM.+KABI<A[gMCca.Z(8:@=7MLJ185YJ9J-4G(^W7=&gP>
1?K5YcE;^YW-JfRZK];02\M._6c\G#<?&-J:9=>5GYcW5d37Ab8,1WX-5O8Z^PO/
INHT4&>(D_=JS8=ARSKAXKb8@\MYNSbT[1HC&Wa0>D:H.Leb4@=dc[g,VIF&3^L.
+CBFc[#fadWS1:H-ZOT_IY^YF6K^cXJUOY\Q;LJ[aSBB+VSTQ)L)Z@A0Qc+PK-J6
5Y^[@AHAc&C)UfbJ#,)PF(NV?N1H0:eLa1bS=A7SMeH8U]]/A=AF,^I/77W</].5
//#)e@>M;@JUW(5XC<T&ZFS4]SK;7g<.L;+Ef@,TF&YfeCB+S=<Ac)@/;HI-MX4Y
1afLM&F(PJ,MV>F9\QLJN+&8#a0LB:9::<\(c,5)cR^J&+CSIX[=3eaT[bd=<?)B
TH]4a4a.6)KgO=UFJEZ8be9adNS,<8dL^\b?=)H0<OL/cTLXH&R^<T^1CD>T?UXe
WRT9^U<CG34YQ674a5O>4a2(,P>J2)\O&fHgBaV-5f-),4VfV)a<&^)O3B.O6;dA
9O8SMKH=eP,8.91V86<cDA@RR)E7-_H3a[VTK+=X(PECUDWN+A5WR7PJ2c28HQBU
F^[+R[8&07^]T(,2IBW+298a3?QJMb49;1E8[RbU=2E?S)E@8<.CL:Fag9)MWc.1
Nd:a4KLY/[?NMN#.&(@CI,9++d>I2LF]MU;TLT@Bb^+3U\LO5HF6gHe2;],56(D:
U5G+OSb9&D-V36aa\;W#aPbQ^B\#?[Z;Yb)M91:#,dLc@;_EDT4V&_4Q=K?6Wg1+
=D]+;LQ_c#f,T?;VC#0Kc_PINV#7[#G^\+7W-&OcV;9[EI8ARaaM6/E,c>W:_<Z/
cA_CcOT^ff+;RTMD8,RL]5JZ)E,e-FU5A4CX9>@6cW2].;E11GBb1e?We6<GTHa.
/]2D?\KMC0d\>3^)97ONGG?e@KBCPPVT:LFEO(Y\VW+SC1X^/VQd+X]MLD@/CZ,&
?fGX1QRC(8DXC])Y7O2(TaG6<\:^O0C_cCD/f7G^D-HRbMGeKR-+O-10BL_eQ6A2
CBJTK<:GY?41MMc_Ka00/L<X?cJS;-WY3]=@6Z<c3)e_Ic;DV555a+d]LZ?^BJL-
8023CZd]5fCUKU56>^e[:S7a9KJ1R-TCB2cPAJQ4-:K]dZ&\W2KgAUf?-=Y-DZK3
F-J3V2=R?=Me/AbO.5+-L=NeU>S8?aEKf]@TSb6B>B;]-cOU7/&E?f.WY[gOTT8a
P2+_:2:/d]e)]^Pb]0VP-Nd1UB([[3^d_SHa:BCN9XU<[(Q##,?08f_F+;=@0>-6
g3cLTTNUR,M5574.FX(EPJc]4XF]CC]f3]LS^aF4K;DcI3e3/&0OE(cNW>WKCTWF
A0^F7gM1YYYK[_68)Z>_4U<P.eR@..PB?BUKE[0+cM6>BX.T/E=XEgLDNeP6P2K1
JQ08R?ODe/IPL>57^M:_OKZCS/cGJL4=,V-eXO<<fY5gU1>B7Q0F08^^,-/HJEA,
R&eQ@FFb3Q?.B.gK3>e9d_[9].4&S/EBd-W_2&F:(S-C.a2M/AWND0F^/@5ZdXf8
@V+UBS)YL@G?079RO/)XM:CgU,T1ZdDc&4EM14Cf;#ET(-<VFP)L/&R6388aPI18
C,+A#9-6d(b=8>Xb,QAFC,agd+VC5N\1QKG-1H)_&;6)T=D];SS]]5KQ,FNJ:W(H
M7S0L,^W.#W2[P7PFe\G[PXPX5D)^f=PH=NM1fIP=f[)P41)P\A9,-EE.WE?f7(,
,g6>c.9+U4NaIE+XDMS&N1e4dO1H+4L+/@+J8/\-55fa)I7OS5VXU8L(VNI<&1,V
A1<93e+,G]e#IafFO)D_K<8gd7VSTYLRMVd\SQ/_?MUa.#DA#L;0b(?E3_Ud5g.R
>;)_ff]Z_DKO,SRgf&3<W==XQ;AQLVD>bC;4&)_bN<Fe2L(KaZD(__1G&Bc;eP(G
XZ2J(d+L@<CJLJScGQ)I?PJM?:LXXC)V2f(99#fX]J[K(.P+MS25I#\L#C\FN16,
Z:EDV<&]1/\E&@TfMT3aDT&e93KDH9\I@:PRe)]c;gQ9J[HcF.FJ[KQPMH^D43O_
c6g2&/B2EU[_4PM5HZ>2G.=&70FQ?9aI00^9V4;e:@NWWe/>dEFNRcY)Zc[d7&VV
Y0YfdS=e,&(a?gTa&WM&=.#a[<RYdd37DHP/,E8INRRS-UZcNW[J?]/L9R/)1HB@
@F_&Q8SB+WP-7G;[\QL&C9GW_5R.K@(3[[)LCR3@B,5g-1[8V3._]#a6O:#M\]Wf
G:3>FA8WCE;c^X/E1BB6?aEK4B_ZA_]Y,_\S+9W)]Ag1Z4OV\@)>\^\QeWB/gJBI
T;FbG##XO;8N#T70ZEAZS9@17AfO4)\(RN>)Idf9cI871_b8=Dg;g-_Y]4([cf22
[.9@\&\/V_UW3>^1Qc,HPQZ<;L5U3?M4+.]-bPD)W1?<P]FgI0HQSJ\.=YI(0GPT
dS#;PV?1ccfEBKAZAH[N[=eC/ead:Y5,/UNa@IgPc]K+9gN+McY7/BR3MBUIKX>?
B=KDKJK,G/fND2]C>^:S^,:.-a(Z2&3&<+f\O^+BE+,Ye+])d]3I68#aYOS(\8LX
AP;>;gA6:cU=gGYcM:BJ,KbP&Pf6X5//3\3#FKJgEW-DR2JF8T\b/WHQSg.AR/Z1
<dbC/#B2]A=+F5XLFQd\QAIH[0T1U]([ZAM2a0abQc,.^fU,R5MOF,gL;(c2X;gJ
e5O<QNa@2/_0W>1f4Y&B_.DILYUNa9fP&DP@E;,aC,W=)e>CWQIP\\T+NMDN>7@g
UDUH5;,AC^IJ2dED[M+<T3KGALT\VKPFLCDFQ[5U]O]gcWa.>GLQ=&<PUY=@>Ub9
B/3YBRe#If-7&TXY74VPX6He#)H/HcY7R?Q:#=gN\3XVK=Ua./DG7C-Hb0cL(GMH
;3-RBGPaN30<V^>9KFCbXc/W,HTX)a)I?a7@YK[OU5Z8U&b)M].>Af\@YL1\46\&
A,JQ+d?&5EEHcP:TYE]U)NE7NZbEF8OeH,^&8R;+Q6AX:-:TD<I;c9P5e_CVH155
[=>F@S=C=UKAc0NB@:7^M.QNA-e[=),9T.+P0@gD;_>TBN;V]M1aRHJfc9CX:?eI
38EL]aA^Y_B3]6(R9>\Je]EG525e7<YaEZYa5]A.a>c&cJ>g6_aE84e,DJHHUg-N
,,-:)[IbS=Y-S@LF?IgQ6/@0G573C.5HGLHa8J3#B@@@@\FF)BX@eOTRL]^7L;c]
:]^35TU:F[;JC^#bATE>cYA8Q1\IJ=;4,6(^/U+4GHV1PJOPJA#,B^]AO+:^RF-8
]W=<2J60^fW>A]8U)+P?eYT6[=0R2Qa/d/K0VV[VdP#<2b5S6;UXLJLYN]9ec4)g
SX?ZU;;gH6/=M920ee>PQ;5:ZLBQ/LOSTIUJP?GRS+,XWK\\4gYM=He\LL2.MVCS
NJZ^Bf:M&Sa-2HB+eC[9<+N)X@D2MBXDP7GL72FHg//1:2[O5EI5W&0BCC17d-;B
#cZR_9a-V:9H2c7(CXcZ+U-E91HK@;\eEKW[LEC^6=Rg;9g:DMZ7)/ORF+e#0eXQ
(0C@3+VaeDPebNXNC[Qf(2NU].1&K6MO;Y)Q0>?J.VI66)\Q\DMQ#,MYLaI81C7-
K/b+V3T,28--3:U\@c<J:,NL>^cDG[[M;DIHM#fTVXT4X[^gL<YK+0GEe&?eD.-X
GcSVC3aD+G_5I+_G)-J(ELBe=IH)RA[MZ,e+R(87;[=IM(>H3B7Q1JDOX)C\LH,,
>(&9VK,H.2]+6]&4^5fGJ9D0:.Ag>Ta]/c=YZ=71JXEQT>_IfaLG,+4YZ#:5/,?Z
91E0<VA@6>a\R&B;3cVH-BOb@MI4<C)A;)Qdb[47(f-D7f<]U51]UeN4F1VD5,Q)
SX6Be&2aLeeGB]^,5POY0_4..==XT3eUI=Y0<:1Qg5@N@_+P-1(=(DAHb#BHWF9K
^XAd#cd86]BH7DTRG-?#a2&Ie5_7EIcYg(]cUHZeXP8NU7+QbG_?a&LQbIC^,1\e
6?,9TbI\8[X6R4dC=cZUedBGSHYQWf0@Q(H+M#9<J=F-XARgRdJb^/+Gcd2I>R@Z
S@N3SCNR3C#DZ-@)=)L(LFC>D9gc49M<egW(9;(<)>\M;dJY^TJ[MTISS_&CN(0P
?()H0BQc-(9.OW3L96,b=<_5W-0T653cd9c^23H/&PMZO/:<F0C\8>VQM_0/fIab
,FHT<A::N&^+?R4SUbfWD@NYAN_<A1ag(=3/HW@a/82P)S+3H9#4>J#[a>BEUM9#
4KbJ[+=D7SbG[IPW9\fJ?_M<dA5B5aJ4,X(V1XPfX5Fe_<A+XPP2K49f;aSAC,@a
G[D\@4\O&c<<8XD3S>0&b.7XB>R?>3[Y674ENR/<GMGbK>JHBCd=6_/YX)463^_b
VeKS\)JTR:P-FWfO(<GR]dB&?[5[.ITC@MRTf3G&YPQ,<0X=.[=IB^](D^K5Ha^Z
)DK0_&2)AW_d\7Y>Fa9GW^9B[^\[.7[ERF.:dM9dAe(fRO1];,g<\47^>;UMS;@0
KO)RKdEK2>^^GDW&+eB:cH0)7M\E7eW-gI_Z>GP3]T=4.YFQ]/0]Ye4;+@5T0>Af
CY&\\g(K+NXUcQ<Aa7bXVf;;ReKEV-+(;b5M-/a@Wg8e]\C?=XI/7bI=bB<B8^Q?
7GP(EY)S-UbV0P58^:Q]M=U:1Ta9;dBA:T;eF73T06-]NF1?]BdU(5.EZSVCYeN4
fMV_=5+A@(0^&ESX?-=&YATXR6>>C:f5fUJ5XK<bK;K=fTLKS5P1OOdD]OHFV@Nd
)\-IMcNKAG_<=^Z<Q53f62AU?_IgD(I+P,5YC33U\e:,IRP5-P;#QCL5PbS+FQ<#
>V5NRH)S25YC9C[2_b2PHWbLIKSGO.,(T8XTT1;\YbbDa\HM)8E[QLD43A]VNOV3
GJVH6>dRc;V@B8/&^HE;GJBIYA5(F)aM=QQZANJ[&)dLPEAfCS9#2JLF]D4NZ4A[
g9Q107BPHY=^cKPDTTXG7+7U^GS:;<g^dTWG-27c#<V1_[KWc4MgQ4@+BR_1:CBD
^fFU2PJRI20R;b4E>#Y=g2QV7((63S-;)ELFMWZF^26\O303/TWA,PYA7\9G&&PG
AA?fIDJ]1I9B3eLeY4fX=(a.VLFgHf2W40H-838K-64UB+C+UV=).IHOU<06KH0L
#1=Zb=-HE)S>>MJdCAIb&5;--3OPTAE#YTQAMG-85(K2b,aXSP=HU7Xa]e__12U3
fPD3Z-<#)VE\NAB1Y[a#0]1Q56_B&ASa=B\3IO8JgHZ^>EdC&84W#@K,82>,8I7/
@(X+PFZU=24UW(8^DA)e/3c67:/UH_>2^J(-V84K;T_Ca]3)8F3SH-eAR\.B.6GZ
1U]LR39&WIY0,L]&E:B+8Nd3AcBGW&2BR\bJ\.0\4:6^bcB]g[L-=5d9bTQBJ9)c
+[W5UPJT624Z?)/Z>a&7^XTHH(a:c=-8CI5R&JJSM&GD996-^CMQN)3/@AK:]WdX
gaTFDLWcHbJ1aC:D9_F]0#P=g113:QR6EaU04.S]3ddc5Y\0GWDEMZ?Qf,O;<+(F
e?(1)-.&X.]SMG_EZdCD&d?N=\;1^]PAIDgEJH(Ye.O@#]5YJTP1BaGX(8/FO^M]
SBg?1MJRY;>88+&:Y)GC6@0eceB>_>S_5DE>9R(/28I))9=@CfgZDI>D26g==BX/
/#a\-:e;M<WOb;L17gL=Y71eaK@50^#DOQG:.N^EO2cI.ZH<I85CeV.1NLd^\)e\
<a@[La&:@9a:ZYZ[T)5Wb&6dL(T-VNT4DcJ(fYFEXU=B.XN8FWJU-V16O<LWYgIK
XG29?3[aY,UT8g9<eO[&ZI@Z)+[M>Sd7[b8^MSgC(HOWKf/CECV8MA/EY6I5C=&K
-N9^\,4K6aUff)+gO:JJ8f0SQ&T=W=dJU.ILW.CG5&\5BbQ8\KYdJb#;fZ]I)e/(
MZ)B75X[^P3&N?Gg;?_f91=_ad=0a1[46+HUYY\]\@W^<QH#.]8f^eUW.UXDC#Ve
8YE/R&.4BfYE5N(NGE[R?+[=:Cc0GZ_-D6?IGV<f[]&4S55If35,-)+cW2S9@FWY
_[G?HR:[bQ(,Zc7@@O-TBGV:eb0/VR88H:&HgGa#<1W;R./&Wa^+dV9E7aB?AEI0
39>V8U=<Q3]W4F<G=>gJ6/b?-<8>Xe#-,[>#d8[DVC^Gd+7@gB.N5Y5\-&gcbdY8
?#<\3.A2=/_FC;aW<<_U7Z47bKL@d,NQRA[<5g60D1GQd/cN>JF3Q#PLC<?)0;d3
2,1VfBdM0LA5:)V--bY#,P.6:NAS#Z3.:?#KeTUJMTKKRc<M+f,.;LbM2@+ZJN(_
=P8dKA3-,&LIV:KI+1N5.JQR;Hf,KJP9JcSZdZgM74.Ne9a/fY)90g<,:4MC6)gK
WSA7O,ZFWD<&.M:(^;bXP&RKeJHE0)dWb]3N-:AS]G0XV2UZ,>A8bQ4B]RN>O1/A
D>e?J))76;WS9bE^9^3,0?;,8W(D0g=;&Q\X:MO^)XOYSe[#:K3X))P3Q@@?@,)F
]F?,S@b/MH]+0CFX0R30(R7D8YCb=:W<&NgZW3>^acgZR(#LG4+C6&=7\]<QD])T
+D7d6eV2FFdf(O(1H0aE.3?bb0^KP<BX=IZb7;.b</OKGcYR]0Zg,Ie;^DQgb2cd
+N^Ad<g<00X@@S_+gNb5I7EEK1KHc821JIb;TF9WA2P7QG&:Z#.=fLW43,I-SNf6
X7XI,a:\b<9]3@IJAJQ3.d#K^GHC][Q@a:AD@\b;T>AM.N1DI^Q\T\)K>4EE)aDJ
ANL;N9YcT/?bR6XVZdHKd&7+^KS((8<>H/V,>H2\6??&d&G[09\R3C.^FC.A_4<<
ZUfYB&WY#e7A\ZV>O<Q7_3QMW[&KV,dUWOO2P2Z.g)VI@HKSIR^EXI(/&-D6Sb:a
2?LMcWRdX39@,72^^@5=DLO7;4Eg6O>0WOTfI@9[^LI)a8B((0R13&KR2f0((G0C
Jg[b/.Q\e1eaeVa+e\<[7E6dM9I;RP=Ac_=Y_HZ6Y217@85QF,3G8,PUfG(L<T>7
81QcDfN.CBHD(G(#.A0?X+[J()9=a@997bHIZ;>P3KgeVU.fLe)#>PKdVc036/CO
(L)4?_;OJeUeE7?<HDe7GXJMTc@THW3Y]e2B-eOL7PBC9cXE]P72a6.^F=6>NG&M
CUDIL^3LX_Ma;M9,:U2f+:7/<SJE\1XX^OEYW)]W3Y+:HOO8W.2M,K>Z@?@1LW+/
.a7XX1C:/XCH&+f.:)Rf>YeXCWE#&gDBeJ7M4KeLF8Wg\L=FJ#<,Rc4[d+cNd[0@
;dYZ\KcVL1D;SJbI#;FM<d9GS0Cg6OTE5=&f8-VK(0e=32BZ3J:XeHM<7^B=[KcY
[OfV>;;OKS111M],A]86U^-0NSPfQH2QAFKX:3)42,E8#G+FQ?Zd=5K]^OG1PN_5
(ee.CIVEHH]MII9.f^]d4@1TVdDTOa]7M:cALJOJM2\CB3dBCA_Q)7Q7[2.4Da\B
3a;W89>B1EKbKZ4I-E4=6@?NC#95<I8Yafb<DPR3egSeDP96O9OU#[gC[DQX(bUR
KB6&5f)e9B3P-b\)\26]T6A,WQ#d;cRWU6FYFN:M_U8b;4#/+FJCA]7:W[DVAK13
b,.SKW@Ec(K7RdD.0T<@^f)Tb]QO[?IWROG4@MDQT-c2B#c(A^KL1b4F&O31]5FN
SUJN+WcRG3A4+U&#cFHWb&0#;2DIB5Q(SHIOOL@agF?MK;4-O^(73DZ91MEQY\GL
c3F6TD[<bXIUQ4OZC<;(YB1f.@8,KEQf]@.(QIEX.0ODURe14:0O=,a0?O8T<4?H
8HbZCgZHD/B6N(U\f@#,#V9_M939+4\3QJ(TT?QP.Q2(SDXGAU,T1-F8>/OQ@=@\
2DVQ;QEf1ARZbM9_g/O+GN5.6MCeDd6IN@Ic\#F?<(HJMH7:XL..05a_L37[Zgf#
\TJ7X>=O4.ac#Y8(^V-5DA0N^W.OY:\[bAH/=WeJQ4Wc8#MSbH947X\NN#/Q93XI
7-bM)&V>4?V2_cdDH4TEYHVM<52D:>d3Z;KHX=NQ(:@I>L;d&3.gZYO^_,DGMO9f
+6+O9?e8;0S]@9K])H8^B>,bFeLeA9ITEU?fG3@RSC0Ha6D6?;IQ0]aRgZ1&OLDA
DR./;W(N_6IA<G^,7FJRX9.dX-\Zb+Q-)KT)_D,6/P_4bLLf<G82,_/P8&5JI6=E
+^I/77d?:+KI/62)+XbT7-_fNfd6S2b3KM:28RF^P6eY/@22+V?GfWJNDHC<;e><
#WL1&@YZ-7E6&&YAKL6DZ]6C;LKcO>RD7eHM,,=J;_U<+#4:R?IBE+X3F7[YA^];
;NKXB4L3dI^SLGJ:73TJ)&?@YZg6;)YUTF?CQ7Eb.K6O8^_710F9[J(;GVfEGGFe
Q\#NN55DDMb)c[GK-\a[Y__UQ/beBB)EfC418eCFc9-=X3a9BK-DIfTCfQ23<XM-
FBM<RBIVK0LAf3K?c0&Y\^3NUIe1D[V4IT-C>[,:6/B]N?>XTd8QZZ(gEZ=1ROTU
ALXZFfV#DI(TAJH?=(AHC<FPSb0,d.)V(2^C=_U#eGUQ0F@KF@3:I&fWA+bA:cR_
fB)8a1;T5:SF<-/RLRWW=3>(KAD1:B.F@\5R.5NHQFIK=LO,_V3;41A+SSZTdV6/
+77Z0&b#A=(e5[eW,4&8V,XG.e_B0Lf9@KPOEB_V3CL4L&>XDKBgbdIA5\@+6dO>
=5:]:>.5,MK6)3B0TQM^:<,X7I]EHP=)^:,\4^;<Z7^eA/d,6[4WHZS,K4/E?LR;
1VgZ=SHP\LfI)8^MPILI&Kd(\C/16KMfc5=&J4e(MAg3(5&\,+adB<#eEAdU[O^Q
B=e7C;6:dP.,,6Yf,241?;^>bPFcdJgVbG_)-UA\:-H;e<,Z[TaIA&).WWA9J1J=
:d#I:,E1&#aN]&_32(2-XM+5e^A,YC@,K[f+Q8VKD;(OMZFaH0La)]^G8_@DALR:
LV>M?eJD@g,fM)[+\3F+D?)Qf6F>VfeaG6\Z.W0eIF,61@>XAf);\=CWV&,A@Ra8
b9e3/NA9S^[-=GFHfc^5]7#:46dMW\+LcP/NBB,/O#_7YK/MJaX<YBL#;YG]Va9g
a&1H/g.Q4YX&C.D=Q4=5_,KC0EDLc>>?;?:CUKS)aW0&1++aPJGD-,\8DWTS^/X>
f@(X91NMMYJ]7>(X@TZI;M_4\ePPY:NVf\CXd[>==Pg&.e1KTWfKH:_ZWQM-7TV2
:HCJH5?Da#eV(,D4=4N&b,fOOM)4V9B8&E2IU(SM3e)f92#c]>JNK)DU95N9W&TN
TY5\eM;@7aGKd9-eHQI^WY\-)3?S4Q7R@8LFRZ@8QdCDJ]5QD@TFI<8;YY&7>eWV
6Wd>:),H_Y+NPY@NUE/B3EdfVHK#+Z(4)Wd9UF^Ob8ULA#GRMScJCS7;=V/L0^;B
-4<?1D.<(d^7]03QgC<-H:UY8X;/XG&)._H[VW:>aTK7-PHY^3bXU;>YggPJF52O
M=H\WM[CP[g2J+c#2a@fd=DJ4FRR?Rf)J)ES5H#gMP)9fSY:(SVWdRVM2MZGKW;W
G6)gJAS:#Y6>UP6<Y54?==B=>HGD)E8g<F@POBRLRcW\HUB<(5V7\Z?g_;@GY5N>
dSP7Kf?4^0OO3H91#f?4C:C<[O@^,a#UPcFK=),CH_O,)E[d_fgO99A9K(SW?[0@
58(Y?a+LNA@V9.(9Y<<=MM^_[<S8VR;79UN7-)=NW##VS)a2DN5\(UJK=RZ7WD)5
N3\f)M:e+cbG_c4X>&KQ1Q]^\Rd+>@.LS:?WT6M;82BC/eZ>XBeb=:0Y(SH)#(T_
UFQWUG=gb6\/W/f:N[/;27:.8INLUgWLHG04)UYT;@(a:Q;>9_OcRRWC3YK<KWAF
bc]?e-Ec18B+9e-8A>Q-dGb:U(+^0a[@.B(,4SccO7de5?ULeLM0DQ3239\F,O1R
Q@\/S]I-eK[Wf5<8=7_Nd[?fdOR6;6;>BB\D[R(I8SA5<GEa=MVF?3fHGIAbR:0^
aUF.K=RI22U\Eg.@8@<B/D5[YJEe9105A&eY610C2RDB?AQJOgC.FL#+WEbU0V#,
<L(FT@#79<EJQCU+\=T+<F>/F]HDK@&ES&eR674Le8Z/92Y]7NC#1:@a]]4,^.-7
E43?ce3dT/SZOBFH/00Y8=g0B7RBK/ca&F0IYM&a9UQ;-)2^NQ]-?^,L3_&IW3ET
8.[IgCcL(]RS2PXf?;L+Z,932Cfc?H/JF.R)419LE95?9>MRHbKRVX3N>COGAD?R
aX,P;@]LVP+#7P\@HW2[f,fYP@Y.0VSc:((I_6T4.=[cJMQ1PKFHV2-Q/@UdE&(2
fa2CM>VUc1]d/HR&3E,-ZF-+^Q9)a8^I-&:IY&.PC^/daJ8]PGc.0#I&XJBdTbFe
G>B2L.[Z0RA3W2YgG3C=FC0<N]R?0WQ[09Fd>FCb8DAM(W62\=S3^T@0@IeE1B@O
Gb/;H7&W=P1(?aMTFJ#+_5ec^(<247a\,\VZNe_ZEaU3.5IT<,\A5LL_2]<CGMb]
S.&5W9WP\^1U83.]E)O<2IE?dg99W+e(2.dX[;cR?\X/bZR0QfU08QS,+LgBC^PE
.b\XG;cP[K,=_ID7A48>JXV=VMd/@0MdWX.bAEF#H\b9,.Of+RZ@0bFBDI\)9.G<
Nb412-2]YO&F=LRa))\aG=X5Qc^/UQ<3<6DR&BSBO>5XYDB\c,AQ6MgF<SB8LT1f
72Gc-<=;aUQ.dO?2,RS]d8U:J.LA\5:/:+P^fH=)a-U@_R2R[+QH^P+d:R393UQH
gY;9LUXW.G<YD5U5N?3V0e3=W[@DM\[+>+;Y&+Jb_LUAA:/-<^WI.f)B;IVZ;cbc
\EP9B=f\>MV?RK<8HMAQJA8J6:#2a>S07D4GA\#(^.]#b;3Rd/U6<AP6.Kba73?S
>U#WQcZY#.YC<K0C?5AbM4+HC=JC??Va67S^H\@-K.g]L]5Qf6T=OFI+HOS?9@/R
JLDGL&5Z\V2W>;-3TcUG47+Yb2X1ceT^@^YgG)F#8ZJb=L)(02Q+F[J3BU(VFST:
b\&S69)84UU_&=\7.SKXA55UPcLMZ4=d0&9SMCW=YML-PYNT=e/Y.0BW:7R[aPa?
bB;OG8/@(&aT54N-U8:+5\#;8J7>5+?6/9ZI1#Ge#>4@F\Wa6d)N=XEWHO>H(F#X
X+PMHJCMe&Mb<JF1ccZ6QBN5Y&Hg2b?BFPZ+U,B60;0VJY[)3SS_HFd,e9?OTPZB
^AgXGU[Id6S43SK>He0IC5]5?dQbeBaNFAI]8)CgM3VJ3<RRIYcW_V,#AE&f_&Le
b0MdObJIA<I-+Mf.Gd#bDJS(EH6RYfM:d,4WP&V?/>-fW,8U@.H.T8N\g3g4P?.[
S&37Jgda^_5Sdd19.(3V:K.KHH<I;75QH^-4JSN=IQH7DBA+@)EZU:bW?OEB)dAG
J.Wb:JR+4gUE/\b/Td:WH[_BaM[O_YB,,aGf0V:_^+:)0S6TVa[.XGaT/e:@Yg,\
fRG_Nf<D7TA9ZC\#9gIVKCDC70@1D<BdXVXab3b1NC#PPQcZ\)YL0bG:fOGP@J2W
\EF>\#\@QQbZ4\=,Vd0.?K^\QgH9[?+D;#GB]>B2)J;/UfcHOBc7-2DF5YY[Q\O[
LN81gIeJ-.60V^#G)A3SeZBPeD:SL<A&ggL3>5E81^_adca.OI)U#Y@?#F7bE<6H
+H7C7NAV3ffa[1FWTQ?f@+5Cf;Bf/VD3H+,R/8YX]TUbA;G(>)Z33D@KKDbU=)fV
@=UN/V^)Pa\(QN<Gf^OX4AM?(dWgHaFba._W_<)V/6?(EM]/RLF)8V1M&ca7g_H3
#0OQFOBAYC2Z8,N,7;UdU4I@VV8Tb>NW01TPB^]Y4:P6(C/X;bDXFV0e5<\(aUU6
BCJV?4Z3B?R[A2C3=\]_5)X^c@ZaeIW))PaH;e1SK<^aggSJ]JM:b<.,_Vc][N64
Oe;QVQV66XbN:>]DKUaM6EBKQMIaZKf43F@I7ZYZ,ab[f/(bKQbC]<=L(,Zf70UK
=8T^.=4N]&4\C=]?85_3Z_KEEZ2#_(-Q\5<OT4S&[W42C=dYES]#MSXfg+]NY)MB
9c)-2\R,JQ9=g(G&B2XC3N7bK=V#KVXa-a5+YeWb(daGG92aL&NSC5d(RNg\@9aP
6Y+0@,6f4=ZKZL(PMHU3(@(e?5+5PaA8fB;DI@Y]1[]\/R3&=TQ@#.>AX-]TEV8=
=[[#NN\R&D-DBMI<3Eg-=N-9DK,:=052:TeO5^gc5O1K2_&5Fc5?N@>:;?3eGMF9
-2]L<9^aX^=1]VFM=a6&\:3e]2\2O=(>9WI^Q7YZ#39HeGFd?=L=O6VC[d_+;IEU
[<R>K+[+G:1]F7^O5U<Jb)L#^\IQ3d49#gT;J0+5c:B)1(W(04c;[O9UKMb@W.MD
Ad1ETXM+Y46U/@3)\420CIC>B>Xg4?0gVPVZ(;V.FQ.eT4U6@+P#4DLggHXPK_\a
@GWQRQ.5]?[PV6O:D>+7^/XN(Y5(dUZ(.fOfPQ:2((0SWOIZIV(7a3LLAHWcD/L[
T_;TPCD\6TBLc-R?NHL/9d4>D:YJ.eLIA;Yc^U1&;g&a]0fL>Yc]9>S+7APK/6(Z
.3UH0U17?GN)2bJ(I66+//K@FL97g+A\E9G)I1.3/4V)7=44OM-<LE^BT,^Q&+DB
d:Q)T93@?^8Ag\1K\d.:/T,EG/217UGN9;]:D8C((WQCB=XTQ77C?H_JH+Sb1A-+
;+<YgFWLYOAP4QJNP.-PH0L4(+Q&8<+VK_5_7]cg19aZ0NP/a9B(d^;O,)QVB-&\
=IRPe:9V@e56?_P9IaQFCJ+;M\SJ5#;ONeUc.eS55=F^a8X+aVf&;]:P@27DCYPV
=)C1O.K0fSfa?b>B-8D\\9KA?0f5_DDc8VF/a[;,5.C^QV>BQ8F/<ABe.\<?4:;V
5B^Q.3TEMJ=a37[].++NBc/>VH8?B0_IgVg79:-3,]e&b<0+GC_,G\U_SYbM&:>>
QAV=K&ACMKfDGPQ>?;5WcQfN;UbA[GecKAZ,?50QZ].EH((:-)AT\g[egS^YV7_-
>+CSTI6?>,CWFLNYfNeb/DC3K\UOdM=6aIM<,b]RHgDOf-?JVb,1,>.UGL9ND<\H
O#:/Qe6)S=P4+(4J@4&g7Z,_[U)XM9Q/>N9eOU];C[N;HV^a03&C#+G1B_gCFW[=
\+<7AIgADcb9.M@)KAQ-WISO(;BNFV=HdSg^cF7>-IT9^/D<4Gg()]>g&OFf,7gH
1/YN1S5=;59c.dE)a9_3+8+MVHOfD:RK24b_>A&X28d]>_)@TRc^=B<QDb-(Qd[[
<bQW5=YWETc)Y[@8MVd4JFI0QU^H4\3/a,gFeaFH./@Ug=X]c-S)KS[VXPT#J;77
g;P#Hb/MTO<.&3]7]8;V-,ZQ]+YZ12624S3W.AACZMR4f[(\;5aEf:#DR#T?I=?L
UCQ(?1@T:<<?>ACcg,M>872CY^/E5Q_>+Jg>X9?9=@#R99X<B2]KFgJc^cKU;,4R
-8/2X[.(KV>1CK69I+<ZR8CfGSEY0eQ1J3g[P1Y48-G7Z0V<_e-1DG-a\?U(\?H<
JDTY/KYcgF-@>?M\2+_e.<5J>2:GJf_B]W=0A1gQ&B.dbRZdGEVA8&+2CV;Wg:V@
YCPf@?5-KZ-R-Uc?AZHfTZ15e13?KW6/<S;W0XFa\P_G_03b0(.RBV<U?[ef^OH:
&HG]2f_:0>OU./PB)S2AZ?D,LLd+b)F\ag=J5BYR-#^)Q7]APTWRY)VCf\AEUT_b
K(K,T),>-9G.9)@4:@R07S)U6-(AHeJ1[6+]#VX>O:+]g46SA()/C@);<7_UMgRe
&B89_2(B]@B>F(^M<TCM_cQ#1Gd?gU1@SA,VSGgWN.(7JQDSK/L]LZG,?FQGVbP;
@fYXR?X2\KU#b20=AW;@?B>CE9e/XE1O@-YN<TbU.^\+-0WX4a./b4fGZ728W/(T
4bZON<K[999[C[_ZV7DE96MFJ_#3fN3QFRF>ZZ_SffNfGd#aC0LcA>_E(#XRBc/6
]G3c:LIBe,6cBW.f<=+=Ef1L4.+g,KJ+AAYcAN(6L11[\?cf=a]U+J-4C5b@O:65
9KBY,8R?[<KO[494,D/&Z0e]J-<YKVaG#<LFI(C##[G3:cf(,Ee=BE^5W^/3=PD^
Dcg@UM=X_>HV2RUMRKO5gOF/IKcMcT3JZ4_-;IEaUL_T3gO,7:=<@]M/Q&U6<469
4G&I-N,fBJZ7-_SDJYReN,=9C&&7[S_<a70;,G)c<3Yf77aVdc3(6_g5<g(5SNW1
FgK#+MABT.)aTR)R(:cK];8U6/<8&Fb-)/,IK(Pb&<bd-9A1#&?4dZMLDT8cXQ[,
TK3-5ZR4)OEgQF>/e:0G)5:9cKF_0GI9B60YgX#T(F#FKEXJf.>=>J&]CU>VMaIA
>G1g?E,H_FNI78a&RS:BN5eUL@e(5<\?OEF58_Ja0CVL5ObXXDA\6/d-8=B.eM9X
3RUT,0S^2ZY(>#;+T5.+<W;db\_^)H.=(D]X5)(9[(&McUDbF:?J.DQ-;5ZR8fOS
_/UWIT2d[])LGO2Q:6-XD&-1+#C8Z.c<&P\54Nd9.=ee]VU6f)X2^H.T,R<;C5#Y
=008DK>Q;:I:HgZ/M]N8:BCKKM/<2MeEDg>3bId+.ea7>(c&cf8KN::ULfZUX#eO
0(?Q9X&Nc(;5&g/AFMOd\<MP^RS,bC7=g&2Q1B=_2)V<,-.(Zb5<[2[-4HeTK\X]
[GZ,L_J;EbZ71ZDAXa4LGfaY1J2JUB:.Ba)DDUME_,-5eSX<dFWMQ.WZKbS/4.:_
#KY-2ZS=_:KC6#bUTbAF(KaK[0M3KgJG;AXSeVFbf\+?g\SNYMHE54LW,R#PXCGc
,,>FWP0Wb,_5BZRW_fX[?EeK;68O2:@dcBS3?\2P+/_AU+/d;8[fg-Ie[4=3EI<g
B6+e1/,aX^2V4e_@dB?^=g)Ef,/F\\)X9Z:a\H#,GK\?0>+=4EQI++5DZK-0GAI=
a^HHCC/;,EGO5N=6VLCN.B0K9E36TDABO,7LS-B0U,.WVF6_[:EEUVEVGZ>f[=cL
N6;,GcQCL)C9CW_d@S1UfAJR126&:(OeUEc2e;KI/JX[gY>S]>:8H@P1dNIREZTO
]>PE3)aWbXAS&,--BeDNFY08Lb.KUS7N-ATXD8?G@YX>a.d.g?Q7GB032c\G\COS
E86X)T(TbK-_5f1bFF7-&KD\FVNU?V.>H2WaLHHbR5#W5NQ,2-gB&LeAf@SUQS?R
Q2E;@Lg=3><^G1H92DD8,CTP@1?^-KHKPY0>SR;&38O.FW(T9HTb0>A_adLW:)?L
RK.&+HM^B(b\XWVQ1^K7]_0a84AA#SL#9@_#-g(EPSW>@Q:fOC6/)a.6<N/(#K<7
RH75aM8412NE/DJS4JU.L;A^>(3(F6GWAVVZHA^G-ZTK;GT:OgOO5H4dQ;_B4MDP
gB+5-eH3B>:I.LGcZ@a-+Te@.@QZB0OcW^d6.EIVE(MTfO,Q:I=4AU?bNQQ?C,O_
0QWF(]QW2-WRG^T6XaJ<M=I]&K30BL+B5Q=-8?(8JJWM(fWP2-d]Kbb+9;H@>JI=
+=DDeec(SAe/(2X[@gOLD^0PB2_(\^MZ[2149U_(2XKWM^e2J<EW6=CC(]11Ja#L
WZ+b#dP_c=;YaKeVf40AR@e7XCF^7^CG@9YMd+/@JH=9NJ&E+JOL_73TIVG4\0Z8
bW+Z-9BW2B^FaXC^YRCYf-_>YcZ(g1>BEScCYHU4YT88#Kd=RU]+LLTCJ/g_@,RN
C,U1DcV4a?)AGd)<OJO6#KNQ+JbIA3O-1dPK8f6JHcQPH493ZfQGdbY]a)Dfe@6\
F8V@PM@S1=cX&a-AMgS@E/^2caafD(Sa\5=7dUZ3,PG>O58R&)>-5-D6K[A]?<.Z
Q4#)9YN7L]8(?OS.Z,Vd;[MI&\:>ee/=(9QB>LH&IVMO<5Va9fC5Y=eFRZafJ1gS
-Y3A1TQK0dD#KH>b&5@Z33#7U2LTcIf8Cb3C03UcGEf.Z;_;(:KL@JCg75EZc^Cg
P>\A9X3b3TO#V74J]?d1<U5=<XT9ONWc#A+EaT)gGNcKC7aL\WVP6Z1+S<4AbN+R
UR:/C3?Ze3HN25DZ&KMbL=:=#28N.YL:;^0DOg#?==cWXaa)R;S\_63CQ(-V[XQX
0BW^b39V[IFOJFc2:gD#D8Rb][bOGZ>.15B<-YcUP.1>\d4aYD<X(#3^4S[=H@g@
CJ51&-V(g60E.T0fZYeJHD6]>dGIR/31X;Z,U+18C9REDa5a?,4RZU\:cOW:21P3
]3#]9O]aa9^UG=MF?52MHEW\7,0<H.9-J6QE9]<BJ7BW9C;VFC0):)UOC\B<#+WR
c^,aF4U((W-?98SL8,&7?9U62]1+TU2Q-S,KQeE+F<b)Bb&4aKXbZ=>(Z<3T+6ZK
GI803S\34X1_5HA^JUXV7_G\)a?T83S.](YWYXfU54XP_&Tg_YHP]_/MZc3U(LeK
.3g3dO>V9>>CVga_]^B@#<(d#VW=F9dU_dPF5)S9:JC5Z;X7g<.(S97Ug].4T>X/
KEE:?6Y0>#N<]dTIg3N+_b?[T/NWT6VT?V;/H<[SMIAOR.U5)__&_Mg^-W+>04I;
(J_E>cKN0V4/[5V>+PS4.>U-CC9&RVgXY<:E-=\Wg2+2S\bO#79)5SKW@@3D?772
g#1#L1H^<Wa&T/A5_\7]-IbO^W1GC#d1g-;C+g8NJ8OEG@7:CRL?eG8FZ_-d[>9,
>HF4_K+Y#2MS<;TL34Vc[.&W_Z(>DKE:(\4X>=+7egU6AO\X:HKAA)/?;[UQ71S-
O)>VG>#JVE5F6?I:VHV6DVONO#OWPMg=N6ELT7dBI+?I+JP&dON_M\Jd?aKUWQ20
(>F-<#HKX2<RQ]b5[d4\@Ya:#\dEX:MfYc#BePg?R3#)F8]Wdb<L+6\BPcC^^f3X
#^-B-34(6@8.=eX542^gONI^\6>-_]Z)F>,86)S\AT)Oa,R)LeX._Cc])#f[Da&?
1Q4=E0.5=Se/J&6+_S=(BU)D^MO(I&cG52cbR+7J=E7P8Xc_U4+Oc3+Ze-+\LGCP
R_1PF<L.O/U#D@N3BN.GD3/,6OS#G,KA_.TL,J=_#L\.,-[4,(#[\d\D7O.KQ#-#
[L3:c=c7#XSYa@>&OKCLVKL>),1I<Gg#38J>eD/HLF)X=RZd]UE]]AKQAR1-8>(,
BZ&>IR78AICUAH.bEZQG5e[>A\;\9eeVVP(GfG\U[;ZBIYF5)cb/WCBgcSdZ,K2[
VQGKX2bU9FFM7L-;9g&ca[6U6U<?:^?Id=JI11+-)0WSK=QcR;.)0cG1J,BX.<.;
2]:@N;#D/8R[>.bC(/CJ&CRRE#2<J4D&)9+&V-cf--Y,B.02)[K92LdDYg?@SE<[
V/4D[_B@\HDKDd.-Xd>Y57Z]P4\SLfW30<U#/f6@H4LJWK4ZT&4@g+.5.+)VdB9:
^X&1Y&6BX=(8dPA)X3FMeC[WL:g]ce54.0+X_;U_&28]3S;a(4aVDZU^28O[5]>)
]?L]FO/g9eXQ>Ie+V6:,/]+Va[M.@E@d@Z_R2_&6,@_JN17RH;cX&5/2V(<bQ\Z1
&F\)D/Z.IYVD/Y&2@,1VSMR52=N[1UB:]6J^Af#0/YgFIZP+Cf78b@XE.^681-D0
LG.e.H#?4fE.?M,)N5XSJZHG8LO+&YKD\YdJ^L>58;T/4:6UXePDW?9+6KcNNC=,
F-Ke:44Q?3A:.2g+N+R7dFK]([\ZU>.30H3Ma=LRF+g8H7FA]f9egB-Mf;gZM0gQ
@OH?J]\.EgVJaVb-:R&+-?3?BA]ca6MJ-,fGAVE[:Qc17bM4[A0,I]97:Z?(JgOR
,WX/69N7K4M=46/Oc.,:VQ+5]<WMYOUS,@fe3UQP]#)=LIJ?@12>44HXQ+gOE2WC
SEXS5G?JB:WQ2[9[&9FY/6?D-eb[gVJK&0-@@IAQ5g<-C(BQ:8Ia:dO-\9;aF5_&
HN;6gBbe>OVbf/UWL7S@XLTM9fU6G7?2BF[76d;Y0+gg]f:4>O^+VRX;gE5BVK+>
Ne9E()EBKKXAM+CHb0VaPXPZ,>8WEa,Z&LVb37,/;FY4g+:Y[K&.14+=-04N9R4X
L=<&YBG_Id_76LV^GU?:NLXW.gZUUBC(H-EIH7V:TPF[)[ZEY9bAVS^A8WM@H/[f
HEB\ZRG^9@X??c&J/O_0cH&Z/<I/XeO;b(7AU#^,C)?Y_a,&\?FMOf98FbMF+6]f
:R627D99C,]N6KI>cc;-Ba#LA0-@d1TQ4Y7T.@SUW_0=?b^>fHNB=6NN:X&RgM,W
]3])4dI_\MB-dVIV4ZUJ/fC<7]096E#P..O,>W\3-4:54>;7?QAd2?X]MLC4aZ\F
GPY5<E,.U[E/E&eLff@SSPV&5:35Tg4M@5A)#/BS&&23(26J;5RYOeN3AcZJgK&:
EGE-@12ZdB7O1_59c#\D-2d62b5b:I1\UO]W^^9700P+60B#&U?F<TXd>(NaE65P
;Q/QO&(.E9ffAA^1g._WIR:N+U[-Z:1M_M@ASV>LZO?6ZaR:-ER0eW?Z^0e<DeEO
AW:2WG>//BQ__9MEbM>84IUc=]NVL)+[\4AV]DMCZZ8J[FHTR>5/<JYZR1B4,O0c
-@7F?d=&4[;Z<Ae3P+0]aDe[M@WZU)bM=FD-Ta^3X,DCL/d()YQQ:HU+7a-g]<A1
NV[^07>BAZXbPJ_DbQ4Z:O59BSYEC;+.:4]MX9MAR)Ibd\#]D/L8).8PRGN.aUI:
5\:FJBOa1Cd:L<>#&^A)R@)@4E>J:]X;K.??Q])eS2BBV7g\7WcacKJgIQOM93K=
J)5ETcV8NS>^)PS2d1Z:Z_O:V(^JB?6+aAE5[bfT-8T]dKKd7]=VK4I6HSUA4WN@
36X..&\+BZIUF49;d/I48.VQe;.&CFTJ;(b.Y/V4MNeMVTO,gU]K/X\32Q)HQT9W
LWL#Lg)QLT03S/&a[^FW[.9aR2QHZ&)X=LfPEb/;E:\[LVQ#I=V@I&+01)]d2+12
OO^6[Pg-bK6+&=g.c2aLb:9^a,b+e^-27#JJMT1Y+:<C6\Q[?EJHKRb\E1\DB0Pa
ZbBRHQDAH_\VPRUT3e(9K^2<a8V&Ed7&#E?;[2^2S4625L1(=5V5Hc1^LYFBN(A9
O&-Ea(>1d3g)^4[56LKQ,0(F@TA0(XEC/Kd_>-])8RQBON&>-]##8=-I?fOUG<7>
L2;L?YIL,:UNF5RZBB&FY4G:8JaPTF[GTKDLT];EaWU>;IQU]&gT8@KOdDHKXF)f
9:<-JD5@)&Q(MNQ1c(MP-d9,N-^f3#H(9,aP6KG9+c5,FLB#;2U.M_/02CR3)HKE
BeXXY7W?eg0^?Gf<fXAWeK4eK=eW&^&A6^eHI+U(<^NaE9TS;8gD_6L81UITXcHA
eaGY(JOLK5=LI(,3VgIZ_^V8LZ8S+GSAd-E?G3MN;7f@_(+Y=6<b[2-bJ>8\P4Ic
0337+FRJDTD/:W_2@bMO5S8&FL3NCU?g:V-aHa=8T>JM&a:Mfc\a+=&Jd1C^NL5W
&W4O?:@M#\M3FPGU6U64KbK(#Le)ba#U2<</)]]/2>1-K5G)\&5A-D;=B:>HRV+2
,N<#bEP.BOA=:8#_TX6?UMVZ0O@N#I,/5]DP5G=fTQA97-g8]f^@ZH58V>OM6K1U
3[9D&6FB0-,L^;K5Z@6V.DS+.31Pb>-AKXC&N[\fb]Q-<2e\UI=^@\;A?X&J[#S3
_W[J,&/+I6Xc45ceK6=/X[e:-WZK@][SaI(8+.g0K4@)dN<#XbZY:^d9g0>VV6]W
^4:.7(fDO?>I8IU(_,EeE]I=TUd;^@XWZdH4AT)OHR2BYOcW^_2CbE<13b?M)7SP
NG?&P_F-fSJT<#^1:[)T5;]:E?(&,7^#b1B^QVgH)C=4FB02OgH/\<Y<0)b,T(67
H;ZP>dS,C-DP]9eIffgI#R8P114L^A:BPJW\__+J=b/]517#.19c<-2f(Occ@:Q0
^Y,6=;F+I;^?\Z^eG1>FQ8,J@3K0eV.cAK@3c/#ODV-g]DW0)F+]5.9aJI@TTaZ?
/I#F3\;dDUPcE?Q+BSA.HaT_6SG9K]7+PKO;D&KcL&=5#AAP/BKa\f.eV5P=(&F?
3X)]7;[Z#BaA_2=Zd63=>WT00^?\HDP=IeXMWF]-Z&/387MeX:A&NK8GR,ZW;NO7
M:^_^g&?47X1)=(M&g,C(E?.eQ4@f7K9F33f/;/7<-DaFcJ;Q:8Bg&34-DP+&?65
?M5DX?A,/PFR\\R,McMLVG<9N/RBc06.^W0L[3.KK5]^?Kga1KcOP\19OX>2>DZb
<Z-P/WdbLB1)JN<VCL]5U3G,AHY.T.P-L)0Z]_7:890SL8-e_+][6[#,VfTSc@[:
bMUK:f#&TPYE4WV=3#V>C_Z=a;PD5,[MOURGd1)RTF.IR+P+O&7@H@&LPBPE)#Vb
\dI=DGRC&[3X\RfG(E:?UVHFaAA-A^IH6DK[+0ac1[^[C3fcY[H.g=F+3Y24-^B:
(5NgD=^-(+^WKUYZ[P0D_RLaB+1U,-+UFgCdNSD4=6]b:Z7TU-NE6FR@cJV_]6P3
0NEKbWT^LSCeZ077<bdaHA]6=b]b9cOB:]\/fQg]&R:C2R1#]HFe\5-f@&.[(65;
c=KM-&50DT#CTO2@.2=QN9.:(HNeFLOP?5=H3SN)VR/Sb[YKNLT67.^^#g?(b7&0
d^?IR#?J)GH+;XH&S;NVL;PB@J@_10NC2LTII#ZgPM&\<#8J1Y04NY0OGMI]#L[d
QAW>AfVVb0cJLL,><Jg#,SF.aDc5,-(5_^X><B+UO9>5[g:_U(WDc&G?5<]OYfc,
>MKUASWL_G@GCBSQfJEgO=4N&VZKF6OJQY_F\9MScW808,##JEN;@WR#ce+\-34.
R-O4Pd]SL=BY/^9(>7>1RE.1d\/Mb]=Zd19eP-B,DC031Z,2VJXX55+_[M;+49dU
Bd59^,LREML20^?d7E^SV8c(+A)5a:1AGH(3fITLadA9E=RJTg@Bb[@MYeC/e[1?
1??>3M:\Z\I<?1f6,H93[Q<+V9V2b&P@0?Q7G/B.0KCUJc2-T:8<=T>B;NGc\:W#
FPHGI<S@8c23S=HX9YTAb-HIa,3D<d<^a[)^=>;3=1=0Z\:NNCbY-aaRd<R=>9JI
RB:K4dM(a[X:R(,WZ(D3V1?UOdPMDM#@ZWEM)0-ZYf-IYO.@,[/.PDTHRJA>&@ZR
7G=gV^b/(]KQF,:GYAI2FS6MG=Y[)NSO6NeU10bDF0;XF&aDK(5f7[;)SRJB?af)
&1PSBBHF@?:1WOO,S1V)EZ:Y9/[/]WK:94/?dQ638:@9W=&&=L4),[TK&YF;RPVa
,+Gd[V2#e?XbI]ad\]JeEe6YfJ#@3#Lc14e&[85P71[a@RA8HF+/QDN)GJVY)gRX
UJ.<C>(,g(B@&.=N(00C+\R&T+H+B6Yb2S]+?fc3J^_bZV16fK\X,9L@XLFJ:LEa
PEPg)^cfG<MVEO8=S.IOebLc9,ILg7/cF4BK0fVI0-+7P&].95)-N:>-g1D/e.,T
,>2=:(HBC<+B,JG#HX81TJKC/9.EH@O=/^X#KROL?K=)]V4d]Q<=aCX2fg[,9P8&
Z>@d(YXX1,;,_,/+37@E7e-;N,LMG1aCfe]>=HN:Y5X_N#(WAScYFG;R.9NMb],5
9TN#F.W)(9)):IF6?:OEVd&gcMBL:C0Q7Z/L2KTST6YRd=?P7BU-N39JQN+Q=6H+
\a3NG^DC<3HMeYS@7:]0H_GK]VQZMU#-8Y]1bFAfeYLSRb3<3<g357M?JZ_aSg]4
c4=J65E]YZ<E\d7_7_]:.G-CHKNCEHIGS_.5_0>df@#Yb8C?P^861?H9<faCI>b#
R.;OJ8N9Dg;=3>;PL0AgY=^C[a_A\8/ZQYeb09fN4,3V]W@3MEE]D[8<HLUGfd@U
7LQD6@O-H>SSK2Zc?AY^D39W9E8KX+KVVLR#+e,NbNE+W&QCZR_8I:8RUK9_UPc]
#<UOdR&8fX-13QEET#VC.,6^c3V;&;TV5BM?.71Jb0GW,[/<XYP1_59-XT&GC7L8
28c^S,)&d<bAUEcA@+-d-BPgGYU=0bA(6^^RXHgXC0b)U=;[&.7bSW9R2W4/P?(^
Teb--P^=<)W<+.&DQC\/9.30QO_0YI=Sc[76.bg/MW09g2=7PNZD>\0\/LE@_L?I
B03ZS[fbZ[/:4aKEM_f;:O\3\>XSMZ>:_SbBS)C8,-dc1:P^aU[;fKef::Z651B=
#9>D>_eEYR3ZKdV&RKZH,:5VYK<9+Yc+g_+a]d[[000&T;2Y<EO&4CSQ\1IAX\,&
.DIROQR[:<;5:X76,gVQ(A[3QJW#18WW<#@Bd+BDT4:@2S8GVbTXTW#PR6a]dPOC
?.=H<JbCLeR=Ef-WBdg0&;e_\C?CRc-cO^R).K0+TF1;3MOO69A=La(I_3dIP_I+
.<.<=KI4RZEb&H2CP0#09e5;d2.[OQ8ZS.(-^Z6=e[WE]#1B)VE4Q.?;NDc68/9?
OS=GP]Gb&cLT/2981HY@HFBFD:GB]E:[2SK>M@)>egf@M6QJ/T(c^HaI<5?K/3PH
.d6<e4S_bM=7]dR#)LYa:XAFAUH=F2c=6ML#[Hc?EVC0=gC8?1ba2255cW4?MVge
LFYU3RC9CFe9XZL6F1VTAQ[;5LL5eFGCaV>T_O9>,C<\WAGA<BT1+][^Yb-E?\_(
4P59KQ.UTJ(AdMILIH/G<3_W^@BD5;@]33SSXV&P^UYR[ReeI.HaO9-N_Y^RdF1;
^b1IA<\=P\eS9bWZ/RQ\FbVX^SGI]-e^+@.#1\R3V5;>1J&C,L/DI/J;acBPUS:D
S-&JP+1f)#YD3^g.c]UM&_/f^JE7\0XF\7bS>8LBA,.7AA1KEY][HGXBbK<1S\]N
J=QL3dZNfVM4L7VY,AGg&:^\O@fF)L5<0]..NZ;(.K^;SPO<;X]F:[-.NU9)e3+A
.XQ=S+;O:gIK6)<O_<IC<8e5f66(#FfEN<_D+0E4cH6)PbK)D-#R8+7+_NAMTA+[
]ZQ/WgM_@HW&<,0KMNJ2=a0>#ZWXJM4)b8D=>]-CR^F<K=e/3KRN5GG[ACOg]RWD
>BQ]>d\3[H:=-P^IBfN&+Q@:@-<E<0[:A?^APNa\_I9,=)27fY3A1M2?Wc:C\KU_
#A2e(_H)Z+/;W7H.#9VXWMOaa>[7MHdWBeZ4g]^>3[5;O^A]J]QLfTb,/T:7^_ZS
gO\:G8EV].X2HaREPQ@3ES8&47<Y\BScV9YPDZ.d^W647=KA1DJ/f;6d\]F9Z0E9
dW)JW^75LH<C51;Y[fU&DL1_N461,N69@VR=^Z4P.2<c(H:b37;O9e,^b_Z;>_/^
UX8@Kb:dA.;W<A<>-9=)19I_;.\:OX8LaFPX\(CL71CG18,<aNVfI-23;6B9[RVK
QO#G9Da8EAOEeE+OA9>T0B&c].]Ke>T76:5/)FA13C@9^6>6JA&4Na^?@)[fM&4O
/@4UQ]DYX8/eYNaJY(cH(fdD(A?E7_4]Q-#\\<^87.0PA;Q1@2Jg=d<D]^aAUNM;
L>V+8E^_Jd24feOTM7-:YLeH8B?V(1&J,EW_SRW+MePEY6>He;>UOHIHR\D9<g(0
F_B4>;(aAS;J:DG4Z\<R#V:9)5?@A?e+^VJU@g2?7RU5=@6AFA=_0R5[4F>I]Ce0
;aAV-\/(c10Y7(#fW3/;T@M&F.f0ED3LE=e3UNBa:Q6QbLGX),L0aK5>O\\J]L>F
SROKcQ&SK3^9A&4e::Y8d95GUNc@R6JAXbLKT]E=#-HWGd?YC=3H<W2_a;-\=_/=
=C_2>Oe8LAbKA33K2Tcf4KE@BC/-TUX<f5cc<:VJ#DN8RNI356DYeO]1>G+JX[)[
TW]YIBLT4[E>DK;dD6^]c0CNY>4HFfP&NeFO\T]bQ8OIc2.e792G9@aJ:9\L2cE[
=YJ#RZHGTCLV/1]1fW=]AFPIQ4/bC4L5QP@Y:f7Za[g8+E]<Y?e#<X@/:WA1[/WY
]]KH1NbST28G^Z2LWbT@^/+?9S)E8/2?\gQTFT;>eXIPP\C,>K)[1\.e1;Z#[C_\
,/Mc+93EC,;<\&2,-Vc5;c16e.g85gaT0[Z>V#^LR=8V/A5G//Ra2UD7B?EUX<fG
_UOMT51PYbfCJ;P_ZcFWB[6OgT^^+c\cW=0&_XF:?ZIAP&50NP[/B9QfcF_UDG=^
9A=@>&3>3[&]cZ#TK_990J5A1VML@R5gN0J>[e(QYCW+&EQd<-6SR;(JAFXBT92_
S2ZSV07>QAaHc)9Mc<4dK69SHfH_#gFXaSMe=>ZU&I&?G54LFBDU_G]DB7G7EAdO
]7a.)1\PIO^4,Zf]FJ7]?GUQ^A\b7:\\X-2T6+=Yg80a/:T8>-,9e3aeSD6(OLRL
.YScfO./-A-J^;M,e?GPMaJL13-<ZdT@e[@dP],UX&#g>PP46+DZ@3b&GLf#aI]0
RaE3^]?V;W>_-/,VC-5,)@VacO>X>g:V6;dB:&,4=H<//?O7A)PgfdOaBE@LG>_N
O1@b=YaN82U_#9a,5^T(L+C;7>?&Z#0[/[_@[-f-Z.f(O.b8UdULf+1K@b6].P_H
Wb]72^O+5GO042YC@T-:8)\3@<5MJ]3Pc/2?0D52,H5MAW[dC4T5Fb-1KX6,fbGZ
BAA9;KG<X7)1H8IA^F^3a,T7-409CJQ^AHB/<,N8[G5O-:GP5+00YTZYO7>=/K5)
_GXfM_JNBeXReQM@P=ONWPgX+D_(,\X-BGVV#fca0\6)1W8f&9Y_=+/\/I^+(N81
2[eZ1P1OGJ<JKMB7ME>e&,.VDHH<QL(]=aSAHfgMg/U7]5#RVZ\E6e=?+51=6,4:
D+H1..G<F3(VMHM4)ZD6T69U\K&B)3),PK^J4#)_L3?#aQ_1/;TYMK;Y2](d?/^6
;aBHAVVOQUI>2T-P9)BZU\+b\^&;J).a8fcH3A;#O3?P=7Z=06+F9O_3MOd+CZ;0
C?=1WG[-b&S6S=QX(V:YX5H>52\\GVJVf^)d/18d;EDg]-E_+1Y#KF[DP\Z<P2^.
VO=M:cQYFIEBAKQ[+DQ4N,WVPF;]a.4cZM3_(H8a:SGb[L3K/2JR,PcW+Z4]bbE/
79(/&N-F?]K?cKHG7U>X(J7+V3c5ACWWb1.Eb()Yeg(.bS,SB5d^ZA6QJ-R_KMQc
4R&8_;f>;f&)S,=b.e:Oc>gGH/S?gY8eRXL6L#^X#2U[Y]+I1M67AX>OB?H,F8(E
H&C=_+/)Ff^U<b:4]KbSU:42:HA_/34@&RP=(,P+D7DQMRWg\92?ZGTZZ?_/<&78
L^&.CeBC<+)1E[dg(1=c<^a0^\MK?_#.55^eX78]G+7RG9aVF1+FQZO9(>)RdaS+
-L3@WS--I]-=EX-K20KMd=O,\=@BF^Z/7YSA[5eVVR#ZR=F]N+3>)_gV=KS.GR/9
ZD7;7:)\F,Q>@.0TH8T5MEf[+T[c.1-9FU.bH\BKObZBY.)0)4#]V82/RXbPL&.f
]KRZRT3ObZ2:49:0<cEb:.=@D>b(a>]0692eB]X3^G454-/0eT&C[f,^=BK;K)8W
[Y.RE7N+,]BZ&JYM4Kb-8(1Q1^+;bfP)P(I>:g.[LT\SA\EdTUaXV.S&QI\4O_6,
.68B8HHFENHR9,_2GB?_Je-fV5NRRY81f<&g0,;C87=<;O6#c?HgUE\\@QCJ+9)V
RI96PYP=&R(K\2T4cH>0ff(E]f<0N#[fQITP2H>C&gg6<#CG^C,b0Q@4&fE_(K>U
LQ=SPID..BMcW4?F?+\93(BD.+HR[G7&N?83J()ZI/B2X&^CZ2C45#/@J8WTJ2#@
IOJA.#UGO<OH:3DR+bB=e=dABB+-EK;&gY]:;.6.@SDEXZ0(.f-.aH42;P26?\0/
TZe.[0=;\ITKf/:_:L5\\aAF;RSHg2NU=a<Y]BC@>N\H>Pcfe6+1eNUX7I3<,aTS
\5_0T-;)?OE/G3GcVYS,GfB&2[.VNc,?DFDJ-R4R#PX[#eL=@b-0,C\L[c@f[I,R
Vb#Og5G.Z,<2-Yea6JNEd6Lf]#C\LRG_-GHHPWf,M&UDGecVOEdVe]bX/CB>JDdE
&HUac5g)IHJO4<3(#N;E]E]g^>4fR#&0>F0-S.&,X+--?Y.O,eb)V<&KEAG\R:7#
&V6JN0LUQ&C.8DRF:da87\:2Qf0Kc,2HD7f:.CUB2GUD><D^W71AG71)L,D7Y9YB
6SB;;20_0]J4UL5.PBfcYGM1N(TN65Ma8@,G5IO70W]^IFc3ZE8K)4ZMJNa+K59N
1f4O7U@L?ZFa=;MII6CK816U[X9d,Ae,9YGN/YZZLP&@=)dFG,))D&QbJXf?LaZ)
g@P&6>cA74Ld_UJ#f--1I8YI<T:?SPKKZg9S6W1B9FbaX[/eIJ>fC;_J:M);FgfM
^CWRZ5Wef2<V4+I))8QG57Hg3aGLKS[;^@NC>Wf9]PH4FWV:^R?0Y9Mg954N/IQ#
8/]8OID295T&R=:B443<31b_S_>F2)-IW,MR<#gN]G0W5f51P_KC.;IT\>RJD#)G
Ic)HF\HYa<e^:4413IGJZEWZ(VBfcPKc[2K-Z&9YOV(L8bX-+FbeTb3M8CEdf[53
FcMRTfF6Z9G@]V[2Tg;ZVS^W_]+_Z=I6c[O//ZC19^>N8U\6C^45d=4^ge9J>+=d
1YM\)aZ[5M=W6Xf<<b?;gT2X3#>8]176MQ2PW.B&KAbO5[_<A/a[(ILd?TM&DPR:
6ZQXf:4e9VZ:>b5O,FSAT>We)>BNN-E=R;<9:,)_]R=6CgU>2P0=cf_PK=7WLa]c
SAc=4g6X^=34bVF:/;_@))76?>0OIZJd][dgdMRZYLO@APe]B=+Ub6_TSQ9VO/Ie
&V4d6T-+3MT8@:2?cC1UL>AW_XFcKIY@#;#3:VI:/X#Rb6UGR25OXS<JS&MaA;bG
\^B7#f.@Q<9c>SSBa,,_fb8IL6-B4A0?15#C_V&fC?R5A+2/[)LFRQ68U7SMF^aR
f9P\F+Nf:R@?YHQQ@A>?LHaD)aGJfP)E;](H@ABD^O25SQbWY3XRaR:bEIT:[5D&
aX8(:a4OA_N)W3R]^XZ)?MYd5PU&1Kd:>YGT?<\>_ce<5>1<9ReEBOE?E.V?>:?a
g(<K>JZ0)OgC5^Q43+/#=DQ@?:f-_6&_XI)M]f?5f(?=B&V.e_Z:ZEE4R[6=UR8K
d81>U+[=NHcU2LY6=I&S8R,Ed_KRF3&[Pf3.X1NKgK\CMJ-G^Y85,T6Q3683&gEg
HZa^]Ac-Q+6f:CL\Qcd;1[8FZ?=[6T_NgOQ[GN?-5J2;PK0)<_b>IA4Z\.QJ7/EB
T18Rc^23Bb//594GL-(3,KbX_X^_3?gFK@+_IX-C.A,B@b/#]EEGU[?AKRJ>-c:?
+?Q?KX>cAF8M9cD;P,T\G.(<STfb81BA6>>3Qc<SH6UHP18,<(FgJ&@[]H4R#,0P
L1]LfJ##=CJ?Y2R/N.cQ[))50V()WT>0>:afgZI4f>)a/=56X2BgI/VWLV=#R_TB
.835A4@5?\FK_4^[Bb9H,@;Tf87OK4/Y,E;\9H\.BR9b3Vd&1+O/K@Va71^g25NU
=H;1_W#J<DRD?9F7_\,,W]=/gbZ&Sa+O6^9,JS+XFNKgI&H\JIS.K_WgQP8[G-,L
XfCBZDaA1R4NM0Y=Sc(.PC?2f_<gDY<F8Ha+WOK6I1>&(b#2)UNQbY;GMHPBCGF/
P-J=3V@(G7EG27ee9)4SbCZCHdf7[V[HGPR33BNV4fW^a07>.7+77=P6=AL[[B>)
\WTVD[=4H5P_,6CG&F1g40)&OZeIQ6()Xb^7PD+YYZ(UG15684F@NSPc&>5NVEgX
=9,I:YX7.T>?OC:gPaDY1R;/-7HTA7_/f/@?I#V_7OIe+@SSQL#&]R,)HTI:=<&G
?MUKHbM2@1&gNM3=3fD,Z-\8&BfLRLY7RP)9YK^=&H\g#P#0A9/,GP&X6&g=PE(X
Q,U]J/_NGXC1eaQLAa-Z0_S5SBFANJ;:bf:O.b_UdWG22/8,gTC;D<JO/Q[C0X?>
b2=d?9@2O0CJOAX3RcQAb91#Lf5IPN@]S=H@EMTbQ.?:5f8110@,2[Bf.N5;VJSL
P]QOd-a-32ZIMP=N8^:_5Ia9&#AF(?37PKg59@^TRL6T&^&40ZCGde5]MgUH-?D7
Z9\c/]S9N3ZFO=Ue^CY4B<_Z;ML6A\R2.dfc4R\KBY7WV:Ae<aDPLgg.R=74B+KP
B]8ED8:c?_Sa3#0(82N1-8)OIY;3f./@BSD1TCS[^R]BFNEa#,Q&>;49@@5g4b/;
+3NZR)bMQ9+F\1VG/eK1R^^=9A-ce^Z2/-UE7BYf#IIHe>.;)W1Y-M/4H&-;>HTD
A+ZU]9-)O+^4A_)b1NAe:&9^UU:X(-S2),;;\\A#KEC:CK]QL4LP+TU#Z0;NZZgW
LN+f3a2M-ea9KCQ)]953V2IEQ0NeJ2\]-(),Z._-I4<.FUOKC4Ee(<4VXOCVHNKN
Kc[BBdFa88gKa/GcT3Q(Tb1J[;g,<#+Ae>AW3SM1R&P^MNH8a@MA_GFG)U-I=Ta&
)JPD?O#N(JH\9X@d?K+QG602.E,]J265aH1g5>EO]?P7,<<B,]&AXCBPZaECN\K1
X&FH@GC?K^)EH6S0G\^fH7.:XfN7J\1e\QW#<./2HZT]=?@<d[aaO\?6&;6]9M\C
1Fd_N(.D-Y+YWA=?K>=He,gN16&Z<2X6MV0KRNHb3<JF\SKdNV5^U\K5DU;\>6NG
Q_Q2T)dC_A;NL+V[>F+g66I^-QY<PV_8-.3#>EOP9^Z6X,47\9U&8?1d:[?8=/]V
.#E^B-cYV#cc.:UJP)9J+:9..SCeA),NA(9OMV7O?eT3^&Z=a0K^HH1[V:QNE#F:
O31_-d2.RE+T50)TJ70IeKVQSIA#W-eZg21Z<^V+BPQ/aI8S):@A-M2KQ+;c?_@L
LK\27&S68\=7McbC]B)_f(:L>gW:2.\3R1&^be;[;c6H(U?NDE[2C,H<H@9e+6HS
3,&a[)XRB(L@V]g^SEPb[Y4G?[dZCLFW_d9QP>QW[N=<b2KQ]S(L;60QH@FAL&&I
HP-UG=)27UTTYE:b0T6WAG&6567gdR536+)7\QE7,/[5<:fcPG\CaeW\Z3/:[7#e
UGJ4;aTdY3d:eg/=0U\OOX+23,0,fJcV<>EWRM]9a.APZF=[#c])GH>3:<Kf?g9<
PR3D/C33^1dW3.29WQ(@f[d8cFYPVcMcT35OJ6QS92E@;H^3@8OZ^)^&=(JG@+a:
_LML7XBFe/5L)>=E#S_K8S>A&M.Z95)3JQ<+/BQLc64JA)7?(Z5@EC9U_G1JU_XK
K4HOMaKUA@>X6HD/VCfFLL(S2(SI6X8b68?LEVYT,[BE[;5AgN69f4a-#BSe\&5;
\c?^14@W/B>&,b8?Q\R;\9>-GACUHBf?E^&XM&UE9KPS3=BeFAH,(Z4<+e&-AYC_
f&M7&/Q=?bL;/Hd=WfDDET\P2eNM</[EAPg#572Q4YeU>E]:\B:U&RQ==5OLXM.8
cdXOZ5LS\<ePKfOf=1WJU38>J.6<44K?9(CC?F10GPVH.A.SYW;H+7GYY^-E^=?7
<)D1YS>7-)]S;bR,-R;AbA&-0H(=]X3cCLYQ.6dG90CHX^SG#WN_X:fUM&:BS4B&
5@ZN#1c8XWH4()[P7URbLSEZB2C.O:a;a?V6-49N^gXR+MYKLAAJV4<3.)97:0M?
[>1QJ4@^e,bN,U:CRF+Y3@J]7H/&J587gSCU)[POIMVDf/[S_<59ALc>=G<74)Q?
.>8<YX>g3d9ZNQ5\7<.MY]CfK)eJ=0L=N22(Be#3<A]Oc/P_4f]N\9[c1432CW;6
W^H#6_)64@8-Bf>?eW@X:U>^?FLdL9Q8WCMO6_9cI=Y,FHbfg<TMeT\aYGDJ_,,H
--NV[_V;a821SBAbA1]dd&(1\</JEX>.c>7D4[PG]83HAM[/10X(]I92/eHH<SK@
YAI\+-c&==^5V)JA.F?FM>W(O&VCWX2ebd)7;4H[<I?Z4Od/<4ZCBSX+YGaA@;Sd
.(-==OT?@E[FJ/K=+&&()<F\g,J^KLcBd,W42ZVS]K,._\+[/I_:]0:6=\&RGMDW
(f9PP]/7VBF,3[GbU=,JZgL)bQW+-g9fY&+cH[B\:HLWRIfFe/4:/7&/I5\)-bCI
11Z<.6Qad1JfR3^.=MY1-4(gR7T0Q<QN58=3,EKgB(gVD;D54\0fGQLN.Ld(\RD@
@_61e&8JN(F#>UWWfYTcA^[WUb,bS0N#K=Q9_dHR9Qf#D^XWYBf/<Q)=e#aLOZ,U
[6HBP:FdUZ:Z\&WERNW9+<f>25e/L^c4W;-X)NF9:W6>J8=;BR^G.^I>e73?Z_WY
UDUY;aI_:W6FfF1]>5IV)4BE=,XU67SEE<^e50SQOC7/U=82M/c3D&^b_bfYY_[)
QKW)7\LNPX?#eaCfK_N::d0,c>@aZ\<)4V@)H#?;(aGaY,(T-6(e9baVFIRSf07I
VCRR#?]AdO>RD1-RDf[UO\IOb8UB[FO3B_0_U2d>7HO,a_55H\IG\B<LV>/A](60
De-</60/Q@O#3T]YYS&gBZBef;GOdGZ80X@YG?CF9dRU?:cEL(TEC(cdJ42QR#Nc
_1/56?2G6;IU<d,-\46Jg4?>-MI2c-7:OP#=)[&P)8ZSE-WdH7>BQPT06LY?<T,:
A4.338?Y?PTDEPT/;-@0W.TEVOd)/(;-[I/aKV(3]6(9OX^Cgd3LC9ZN/_0Db(af
#7K]#I\N7&5:A<4<RXbU=X>)^Ue6X__B.^dIV?_@HM_f&FGfDXbT(S[6Q@Pc+QIF
PQW=8J51DFQ(0NC:EF(>B-N=P2I_?#DDM3JKB+)=P8O@:N\(9b)^Ee:QN(3<?;EY
fdQLM7S595J,.Td8R96]Q<+9SJ:X<),#ZNe1KE3XZ[]D?W[&_&^^\Ce#J9a(O9<K
OM[&bZ?g^/_IWc0?#feY<_GEZZ81:2;agdfZ#F@eYMBd?=ZVLTJ^Bbcf&C78PNR+
I7SH;9V#;U5Hb//+\VQgJDE)Ne,3Zg4_]L;-fe,UIV+-LKR/TK[,OgO5>af;>e65
JdPXNGgb[2AJJY[]+U7d-R-1@QLH;#;(aE]D(I^G1]U\K&GB4M[WNNKSgJKLRV[&
.BVa22.RREI&.dG3YBFPeZ,9TfbEA(C#1@L+Z]CdO=;.S?b4HC[I.M?62d<J+AF:
R&#IEPM&/Z-]MC05U5NZ(]g0)RVe&>MZBGUfU\.YU^5Xd_[(9@QR<bP)2RQF2N(5
0\#)D(ZcJ_#ebJ))RZ/UY3@bAZReZ/<.0X_ZG.UVRJI2^Q5QaGKAgQ3/\F(^=LX7
eH4&P9-Z89)CCE9VY.NXT0+)\XT7dg,d,3AJ4YQPE3(QESKC1WFP^#UM\=>g+OW6
EX1OJG,Se97RJ\:PIMQ0aO48\2X>8P?[Mg/03MCa&d/bga/-#134Y8D)bI&R6]U;
6DS/Od=A2EfZ?N7YX]=4SXPT(I-73^JC.aQU6VHa5C6=H&]-Se^MVC^L8TfR@]2H
Ua;08)W328.@0&M7_?JYOJ/Q6O76K;Q^5dXJXF_F:LU_91PZ2M#GF;>1E8;gEaZf
c##K^A8:4AAP_HeOPZ4K;1K4(Z<Y.ZEX^gCaU2Z(,YQV9QCVXS.1N/dQ,cAV[2<.
YV6J.IAc&2;AcT40U7VOXFU7\]2Y9IQ:W^>?SR3c1MO8^,>bTeE\(cSJX;O#]_R.
MQO@2ae]3B8GNMR:bP?(ZLLA,7UgaQSBPaJ>a/\&LW>f-X<eUbZN:#U,6161gbXg
MX7O=,FgeF#eeO[OLGLDf-IN9?Z->/EL[_,^/Ic>+=;[/B\-DIgN7B]#aOE#Va0R
T;4]11gD36e,f.CQQQ<T4Ad9#6>OUeaf#.&>C7b2N>E^#7e1K>cBX/3AEEM-3+5,
#[?K#eZN1#+TP&P10[/_#N6>-LU;/3c&I<5c(.c@_c9^[QHc1]W.(1d>G]B9e#8Z
^DYFHeUbBfcNd3(^c5M(/c-^8_\T^,.AC@DTBL?CC4>NKgY;ZO_/_@Z#ZD=L8()9
4<;G\Z6UZTWeFKD8BA584[3&,M2UDVIBHIfREZ]T:EW@_0WJ3SX>R5N/Q_(3S<+U
WM3/(D<dAc5:\H\:?#b?/cR-cb,KGHa.]RQA#38OId].\A)XcVKV.#ff#^=WTYB3
AKRDeb&:?GR[d=7+H:Icb;)HSS\)TKG6QC,CU#1AX[RUH@V,)>Zc)O=A^4G#T\Gg
+I/[6TO&:U\WR7_R3_8>cHB^Hc1WHdc=_=O<NUbKDMWJZE1JVH:DFOB\M6c-WCX^
eBKWe2\-A2RQ+gY[XZ<OJS3Tfge-=2d>Bf@f\eTR)FA?_;aIL2^Z&H.O.@d;5-3;
PaeNE/7,T4+QE+Yf#H54YQBd=L?OG)c03[cL_.<4ZR-55<JRZ:B-ccRTe8fRFSJR
8[E#MVHdc[>68O:AAG2M32TB85Z/ICWM)d672U/1NIK&46\BG4>-?53&G++JcQ3G
HN:8JXV<:C;-U:THG1eXBUa,a?/_agAD_=@S(YY/f0KUfTXaS]-&U<cGODAD(##c
@A_7[&SP3/0aFf_SFB(DD_?>-,]Z=H7(D-V@BPY-Bf\e;\K3,A5=cCJ4OM88U]+_
YCGESOVZ.Q=D8_dH;LPT4,NRg54dQB=SGXWL17c3EHGRR\U>bT_.#d#fJZ4g^LD>
T50.Y2G)R_a>gQ67O[7HU9d;[E>X[5]=1Xe(#G=5Y7fbY2MFNQ#D33Q6Z5-?BS7?
4PgII/\aYCV&ZG@QOg3Ld(O9=@C9I;TG,ZVS>68(JeTINgXV&\IVGV72UF:_(ALS
BI\4.\Z;F#X3L84OX\@I-\RIgQeC74OaIDf_b<O^F?-G&(^?7L[J48MV55.:SAGU
Tb1DDA)J.R[bA@NK#?&;O]4\)OI#D-1E<)Q33NCBR\GW#76].#H^40N2HFfXLL=S
?;RF3[@WcJd6D.@DR;I=fFHGBVa+g/?6Y58ZP-E8DTL&HR^QEB3_C>FIDU.FA@a>
>Z25APZ]&6X1L;(eE3)XRPfC?Tg^TfDVK,PF(44(H:d)6@,88c]/@IX+eMS:KaF9
M\O&5V=\eQ6L0I49MLFCTU&;&7M->D,6OQ+[E(95_>^C3XI+#AUf6,T#M;2M+e)G
0CG1Z\?^NCfTDXIM_WPV-f@QB:L>3?>?)+,,6Mea2g-F2OgV[6d[Q=;d68VUEdH<
L/??\=B.\UgUQ.4\8<SFVV114OWf2b-B&,&d;YF7]4f=8eC?UL\d40Wb@B&.(FM3
UP<=;U6J&(1MOI@T:VIR&P55LE(7S9BX<..0f(6f2_LF-5ILLG-OD7SeL\VJ/5J>
T82U=:9;Z(S:0JR3JCVWETG>W,YCHQS^LW/HG)a]>@W:#^f.b@LZ=N+fD=U4FO6^
b-B&,CFJ9;WS@H4&ZXdET<SfLJd6<_M4E>bT3Q@(MXa],cDA2;77[:MGMb>Q3..;
#BeD]22SNTWgG:f?035^^H(@af-@KQG8IX:@][cK:-:6YZd=^<WXQK,P@1:GQYbC
HUF>V8HMPVO,#TV)>O<HLM<&b9:cZBJ&MJBXPN.KHEVHEGI>TP1AWDY[,PIU4A0R
[ga+L@g]UFZ-@aWfA)O?GN&;9DUbf5\GT6_I-YJ/:U1_TK[)XFPD&E<LPJ1>Ic9G
11WG@,FD?[7ITg05DQ0.TKUNJG?_10#VW4P2;5]bB88F-(@4U]::gL?>&GP2]30d
1FTZ?HZHK]/=5T:@WdWOYNY)(P?,XYX9Ef@J<MK\_XT]5/e9QND&<DEM)@2[W,(b
Q(-[)c36DcCBcMX4YXO/HG#&^M]#VeUO:E\a<.V0)@L-+;(/ZY3>c4<+<X6.@)^V
>_.HfHVP?8MYf#Ag&/Y@Y?ESSAFF=Q?^-9?_._J)UNW6c=CdO.G5AeZ_[-H1dbcO
RH.A7&;Q,JUXZ)C#@>5+EO>PI/fKK5HCY^+7#)JOU^e7T-Y1^AAAU^eHK>gCS.7G
BC)4#(.JbXXL5+BK/-bVf\\a;7/66JM:.IF?^Gb&[-L]1DB);dB/WZ[Q4L/9<Z0E
4AJaH(M6V_d__1/=5_\^M4FEJKdNKR@DU-\TNS\YIP5/LH)IgHXTD6T\7M65,bX^
HI#&5E,1.QHeYFHCVXc0M_+S+Q93]DU\X&5GEDXN9&UB7,1KSd\2X3:W3A_e9NK(
C??QL0@S0/FHF0W^[#CUD8WFXF\A;/aAN=]c=]g2Y\(C_TA;CDHaJ-(PXKc4BH3L
8+QJU@ZKM5/8^bM>/FLM#IVL@IC-M)5<.\1X[Z8)H-Of+,3gB8(H\gNPF\S&<(NQ
e>\d,0YS[RJR1FY^39S\U7/&^>a0P/4QT.]JY>6^91N/6#AA;?Z2+TC>7&/^2QIO
-Y:H_TG(@F<DK^(>_K9/:HgK<QLNTI3c2WI]U7b>aC;D7HO(:>e/_7X>(<Kc7>K\
gfT4gI9H\9QHfUg4_52N1H&P5/.:+EF9UUIXZ>c/Q#5G620/,&(9Sb#eWMB=CO7R
6/00a0EG^PJXB6d6[5aIQXVZJeYS\@>M&1.+:.6+A-_:SELb?E7\f_\1.EgW[P6U
8Xe)7XAQJ=(.0[^Q+gZb>X5/I.#JCf=FD[WPB\cd:&G9P<3B<@=CfSSWO-]@XW7H
+6&>,_</:>A8eUEP5]eV9\:-Z)9<+]6+a^?=-ENLXU374H@c4Kb,&]70.=>IX:JD
JD\+Yf5UK_Zfg[;?4RBK.[6Y6-gKX09?<X_eWY7?7;1aIK&e[/VE(@K8B6^dYH;]
VH)9MPdXb[Z0#(G849UZ//L]_3Q=\AF4;gE7^:REZb+Vc&T&W=NM<U>]&g@-g2=D
g?W6NTa5ZZT1W=KGFb5J39RJ@7R?RdU\\+BP5^V2I1MV4Tadc)J5>=g\g>?V#/E^
?0>\9;KL63(=f>&2fXAB8.AIc^[[K.fS3O>(^:09Kb,5G_5M]QF7>OeF6^Wf2YeK
1F^_KYZ^/T<UBFDH8+S_)K.]0F_Nf03f?#A5Y5<_L9?HDZQU.ET_EO[K;N7.8C1\
H9VENH[[#K5<f/8NMQX-D7?<(FGFLOQgL&49K,:Of8]RScFaWf,_.a^GL38-#b3B
:a<2fU;DeH2C<Y@-^6;/PEW[EfA;FN?\bP&BZQ#0\9GZS&YQfZ?4fX6KLSWE8-T]
0HKL+IHOX6+Cb.._Cc9ROVL@P]N?V,VQR8W/3Y3WOI0\dPdN)YY<.088L[J_<KE]
e)8&YTc<(SUNDS-+AT,.LQRTHI5A>WT+_MK1dK051;LaaE1N3cR-<[FN7L^MSI5G
E]f&\9,I5W;M?VbPfMd:R=P_9]U@]GIP.QA:eQ#<Y#POUdY:E>>6,I@Vb@/bCE;5
EBX_^2.0JFVH^UP4LX^LE0HG:)f6B_[RCfE-G?PG<A0@VB)U6W<dIIY1HA@9?07a
f]aU0?XYD-6gT]S2KP0J&:JW)[17)5JO9657]BQM3&&LRY)U5G_P&=3cB>&P0;d4
TL<>9SRH3NXN8E(S[HPSB(HYfLMcVAOY_31aHKYBSD:J3GC4DPcC^-[&7]9Z;O<.
&HW_?\@9OE7D3gM40R,[):0d]gG;?UX+6^4;JK:KC&Z8cg8c,0-\f<22fVC8Z0>>
bUUAd.V=P>X).;B8R-1b2N7<]OYP;Tg1YaMRA.7E43C.7g/5]cS15E=8IC0.e,B/
.P5H__Sf39,K/\/BI_TLL[/fL;Kd780T<[QS5a.7H:8G:+[L^Lg?#NcY>4LESE5b
XAN>8e:Ka[]A<\d8?1J<3J#3)McRdTa)4<6H+b+K9agJgH-dP1gWMgbe_#D&&LEG
C[:9E,X_O&fQbOQ8-<)6I5W0_C+>#]9=TdS=Z5UJK&eTZ4?O_IeR5>Ib.F[)Df9L
L#J0,,6CA8S#\5R#Q[cRHG\OM=C&Q#?=&4aY0/TRU/+Tb;g;fEDLA=#eN<KI2&_f
=-LOL.^..-XMeBLMYJJ(8AQLV:Ed42M-RKD02NB/>9g9WYU8COe]Ebbb3<AIE[U>
X@c;\DZ<_ZGD;XFV^H8U1D#bdZ&Z4[HcY3QAE.+1]3>=<LBEd?F__4&39.T@M8.B
1N@NB\,FG.L5&)4RH5O6_O_d9E5a[gC=^O7SPKT&@@T-4^JA&a:#0,F-AP-aM<WU
?XZXH)M40_&A:JEB3,J8-=WaXEBb0YEcTg@YZ)J&E+.H_JX7TdM1(.13;B0@3[37
,]16ZHdT&(]eCf&9A^\b#3ZVV:MY-,MJ?IK59fV,@5M36bE7-:TKX+/D;(c7U]g>
80C7a0T4B_2(>]1R<a<b9U1@3b+>_+e6Gf,(PFG3=M\(M82FK\B?@[4-VI:Ab>^a
+daPfZZ1:5,)S4.HVP95#^\=VGQT8a/7#.c^AeKLSWEABUbCg2eV7HY>0,YeKcg&
fdD&39=A7_<CU3d@1^I>ZT2WDGO;;]8E1T(Q=N)2Uf-5S1A2#AC11>RB]:D5eJAL
?D:A^)R\5O_YORS(+MS?N6SP7T0K_)BRX0@&;B(g9e0UQ=RLJ2EV:JTO=#d7)--[
?M-Fc/?QMO,Xd(9W_0?6aA+0IV7N+:NSIN7Y0Z_+O4#433U,H].0DfJ([:\:c@K]
^bgbXE]Za(+f7e-G#A#UXL3(?MBOK#-,U_2[gX-+BFH:8?/a<\6--Y=S=\J.c&P3
)3>282^II4Q+Y^Q^eU-WK@RY.XMg-W+(QH+TX;C]ZQI?L/@(KE6;(([0T?)9,T>a
PLYHXYM;=JLEM0XIE/);LE\6geXF6&d,b-8a4YL,5QbAU@MA-)VYJM^Aa>d4aac7
TX5cW\G?d?.Z0U?Gc:;7A-KaZF[RB^Le;?KSVVDTTg9=P>C^Q[a0V52If5?IWHgL
b2LC/G@JNCf9L@T27B:^6K=<1=d(c+R2/G^da.=,c@VY([EP)I#UOMd147ZAc\PO
+:fIScC@cUbb216FBU5[0/X/#Jd8U.9Y,>(;V=b2OgYD;5@Pd6,@]Uc:6[Sd<6JX
?E6>E5H?XIf/IH(<4b+YedU\:bD=+IC):gMLWQ)M;Q#[C4RR&,E+aDG\E,OeRRF:
CD[/7fLKTA[1&a&6^JNV+H_OJ_<JH/ebDJB3QNb\b[T_,X-#7@\S1[WX;&eQH/DT
8ANTgWdLIY]GIV(HIUTKYQM-<K]X]c=4FS>aXZ6(d:\Nb&QE5^+?<P^::Fd8<-P:
:M5AQ/:FT1N)_Ke/BZ4,4-/Q(P0F&KP0ELgb@1O6fb&NYZX;<LbH/MeS?ML/Q)bD
##N97Y+GDFEXGA?B1@QM>W:09:aV[3eW@A-+d)&f8Q)7_G:MgTHF.Ib^-T&0[g6b
FbR.^2,:cQf@KY-,U[)[7\\c6^\>[04:g<?5U5e6B88X.]3-CKK#G8(,<.JBI7Ld
aeO8Id>3EcaBff75a7>+66:UJGI:(?YJ0I(Oc^]4ZZ;CA@TK-_:Pd<MV;X]J7d3Q
CcU[cE\Y/1:7D<c33JdDa(28_X3<O;e]N_5=FIcS;@g^))f6L<?3.RG:62H;U<UV
N,8UVW+fOEYWf,]S2=2eK)@)##dIY+9+YcNXf_V^5;Q9)a@\C;N<3a^/,^.T8[/V
e57bD_T5DF?.Xb/2VE?=>DTWD_=YB;a.<Ha<G@e^[^4(d2ZD#)L&@<TT-P>f)=A#
M?>fO(-JdVA,<ZIQa;EP)#6Z<EAG&)Q?U\=9^.H)-C?S&WZR;6ca\gQQNZXOZSfB
EO>[#-]Y)F-I#TK0A]P,XAPO<,SLP\CZ[]Y<MUVRZC\<EdAY],eFg^3Y.JVUEN-U
=.ZH]Yb6/]3Q/9@)/FRVVbg0SMI:9XT@_4IBQUQC_/+eCEaBQ8e7fQZb(Xf33cPf
+QGg38@OU.VNI6JIP8Fb;2AA[WcX\)M0M(OOeL:E0+ZG?0808Y0_\Z1JZB,BVE=)
^L72TGd#N6+>210RGAg,+fc77aBBZ/dJ+:=QL)MXfDVcY[WB1?SWN?GD?[c@8B1]
g:SD>T2JVS>#<f1_\1LJN+J:5TMD=#KJQ9d(>DD[4],K2HBWQ1XT]GfG?PB-K4_b
^RF7<&2#FM1#6@CfK>M:DR6#e,2MA]P^B=_6^TWGGe(-GSZgB^ZA:M]e6Z:U9HFD
;T1cHU=dJYSCJXTCY5/&Yd)IWe_>3[]VFP,_P<5V;ZUUN0#IIgM<gLX^5HUbEfJ(
R>6]X)9\K;8WcA&aL[aDQ@6@/4d7]97,@&D?J2)?Ad,E4:d?RB0U>?0MOd#[W2Df
;E(;bR#7)XWAgZHE;EAfb:+IQgRFQa9Tf(\QFNZ\Z.ea,f07;+?TU7gBZScEDE,7
:0QW83X#OG6NL>a3]\PNaUIF6B_RT&=\]d632Rd&KcVF=)YN1KfJV;[<OD1Sc]Rb
/0@W5D:&0:>@WTF<.HS05^WV:.E#KL8?9KI(2L>f9YIVSC.D1]Q.=2H1B0Y;g\g]
Q1aA(Z\#8Z(_@2^_@5FR4SCcSU:B3)>2R(cd@JZ_5\B0;W:VRU=H)(EN44LO(-I:
1afR):5Y<X=XME,V?M?)H5+1/7a.K#A2-;RfYEe/).(M]29^M(DDO)gTYcg-aB9A
2f/+UOG7>\.E?]]O=5LDEE4@V^;P-Y/S5=L7FKeJ@a+T9cED;UQ=)@4DgG-gZJ-4
)NX&eYaJYEf=W\5HV-744_g07aEY?gZH.A:)#>T,=[M9\W;KKfV\d291L@ENWPDF
87<B-cHg_MAce)X6f=>,DZ/:WFJJX<>\T:TK?1;R^4&(f?dNdMe8@>b,:1ZO3aY>
dYVY=NEb3\-30[;;5POg;1.HEXTJYB/HO,^_H7Hg18HX+2X4:XBNb^:JcDRX4Pa4
=<E5]WX,QC_OYLL&9gIMT0NTXIBd6B/IX33?(&5gVS<R,H0G/A^)G>4@.V1,b,?;
&,\>gL6Y&S28#gdAYTaHAU3QKFJ)-6_]Pa<93+O?,EZc,?-CI4d41NcLX7F#\X#S
Xg=cc[dNY;8Re21@E1E0DQ3^=;\7FI3Y]ga0VCaH_&g#b<G/2+O2(-44(D>9\TQ-
,Iecf2U_Y7T=;;[R\e7M0R7XIIBEg?T)9X&Y>BQ5#=[#-?f=R;T@IV@aKADaY+H)
[02,KKTD<H2IGP,Z+>5GN]\Xb:cD^a2N<A9SX,G\BfBUNI+C0UeJ9R&]O4SJEKL-
LFeGC>LHT_4R>T3E+F<KIFVA<E9YW5TQI4T5)BL04V:W/HUUJPQa4=d@LCa?7LS\
FP36EAG\UFC#\V0/JD&[@8>_X.(@/\>;^--bXT47<BGgPFX-W4.e2</@WL4:;5_S
+]dbf4eUNfEUZY6OR+M_?2ZQ^J6-,)31.)E,.fTH=HfEY)XNCIRK>NDB(Db174_=
26[UQI/Ec\+(0HEJMQHYEK2F_Z)HELN=J@5<O.A+e1Qf-GE0]/<EQgN5#DKW]f3]
XGTBWF4S6WHTd#U8.5YSZL=7NQKH,ZYSRaWZ;XERbcIBb0:G71eNX)J5bSTf8ZUH
Bf?^B6.eDdG66baH9P,YTD3A;X[L+?NbUG?+9.b/IOM8#BKVdef^dPC6dGJ9a9MU
ee<P53>?Re<RSN-F7M^>^9G\M^188-^4.EY,cV(6,VR:dEg>PEK2)cD,VP#0K=WG
83:Q8fMQ?LF]SI=NGNPW\cZbIQ.T<#GO<QQW#\F5[gN210Z\>260JRA-/GWLR]FF
SU_0CeRc>60Oa6D2^H?4bWEOgHVAK+LBY_(#6#U:C;I.KP49G6=9/e@3DAC>bLE<
(efgA\G-O.B=;CP4DC\4J+VSN2U/]SZIK[OQbFWeYF[H#X-e>;aFZM3K7#M/AYGM
<3E2\)7V83;UAU6/JIZF,7,D3,QScUf3B4(bHbR+/DcYPGV\MY]L.?F[G;CZV&ga
P:f_\gKD>JKD+4/T7X1JK0;-UPV_?92LB=f4M>?30@A(@7#.:KNQJe_<PK1f8g.>
D)5.fJZ;Vb-V/F\RZUL=EZ0#5TD&cDF5c\([=TTDJQ2g.A2M_9AaZe),5C><CTf4
\DY].eJLP=;/dbT7ePY+\G&1O1^\6Tb=<4[&Z90@^:06(=]A^.,H)ge5f#WMN,H&
VI[)B6,@RSWAR-cP6+K..DP,_[&\+]0;[YJ(QG7X90A9TIX;F,f&e#d4#Q.;?+&5
]fN0J_8/NL<L,cf+_D#+P6TF56+13S,4eTXNMYH98)Pf#;[YSIY(ZBdb-cfV>b[R
1Y:1O25I0(W/WB[M8CgTA5&)@NA6F<=(.PFg>DX,C(=\+-T+.P9Z0I;C,f;99.gJ
VBKa7:@8C1PYa#>)]DPY5BMST.g)M+d6<+f..R0O,bf4LR3@=R8Yf=5_^Cb.1-H[
+EdXAETYXeN3+cRfMecTcde>02.E&H\S2)9Vc43fUD@LBf=-K:754&@G5X-M@VDB
NEXS:NIC-LQ#OfWU^:b&;bD5_,BB9HQ2Y7@KLUBOPR=FV2G;?WbM7T=&:Z?gA<eb
[cQ8f]LDGMUMCDG]E+__]9;V=<dEIV@a<W#W0WdG)/7ICRaA5]@CS2:WfMM+dWbM
4I+/>0SZHFAaSgT^NBJE9:Y[3F2@SUFD7/?WG/VQ?X+7(9X,?NFF]G=c?+?V004(
-,dXAQMPAc]_0H2&AYa.<B#a<#J:a]F@;ZcM:?^L(,.EacYKO;;Bg(0LD+Ee9GY4
g+P[[?Y<cV1M&YON-ZcgE=.>K]]7(e/RC(PBK=KRb)bd\LA>FLf3ZK@L<[bKJ/g;
O^abUgfM9F(60,gd.aM9^IH0?&Ie67FSC<+QYGDCRT]e7^J,W5GCPEcH.Bb/T(U[
SLW5AD+[/-Dc\FZPUa:Y#0e\(E\Tg^ff+5S8HP^6>B)a36+bZQ,)]XSC]1&P41V]
5eg8e+f^FC@HFUKd[Q)_WN@#]e8Y.BS(1=)]O([TfND#G5E,2RKea^[dbaR3]F4f
)b2-0J=I/89c[SK=Z9&2]\;M1CFCS03K<,/ZU<eCf82TPdc9R-.DIgc]STFC>-Y+
+E=)f#LL6WUJ^M3(<S_?&ZUbH8:]Ga&/VfZN]c@-BBb4M@F_XegZg+_G8Ob5)HdM
:)&=aKU,;cgIaT,86B[;^&S\X809;_/WPI.0C^A3]E620\]3WbVHQT\KVT?GM(44
_Gd,feND^fV6,Uf/<2c2ZWTKXMAP.JK]eM2=ME3AZ3F3G<,c)5\VVUM,\#P\AOKa
NPO7GB\0Nea>Cg)EDU^H3MK4^Pc;G;N]JHA36AM-Pg9&375Y:PB<0YJ&>)>/<UJ3
Y+9?-Jg5TAP@d<CbD85U_<N7<aDR34d/5Fd\>/)e#]TBE;N2QSC#2CKg1XQH&H)\
LM0R2[ZZ2fI+;5O2=@aN;a-FD[J;?d@HFX]TcZPI;RO2Sf605>Q#b1c#?X3:RcZN
2VIG8&4VM9C=Z<:05BG5e3D&SaBI.fJN:;9/AG+77MJAaT.OABga#,,/;:>O#]7e
VN-dPV>K6]Q\J@WE;79G91<M>U_S#bD)fR[(,\6MVJbGG95F(UPKDQ,/H8f],1M<
P0CLNG4:UV7Z;:AT#:)bN^S]CN;:KEO6FF)4,>3+[0=]L_ZR?d.ZM&?Ad[f?C[f[
?fZAdEH9O<TB1[e^eN(6Q-6N&:,5G^NY<2-#Y-P4\\0:[LGff&-OW8@UWJ1.^M3J
J?<gNL?^g:U.,UYH,>9K?\8(:J+PDZc-VKQOEY?ZXSKM<(fR<S)_]?\6(9GN@F(d
9a74OTUOKIe\aUO.gCQab4ST>I.E43U5.c&;)>SBF>-.#UXH]=ME8dg7#M;RKOV=
6W(XB\O_W(=A@C,9+S2:>]dgW(b_^][Hg@A:NXJ7SGL^MUZW=b:1cTJgR,<U@P;T
6aH^,F05SR7P>4?R#-+KU+CXTY/IcZ,B&5Od?2,Y3/K&)[OLJI#MK>\C+PQFc9=2
HZ47.bVc_KcH^)[g9Y5XXPf&1?;)+9e?2#Le8d00\=O84/RU8GE9a;NOBAfC0/-&
[e[a&&=F/X<88:e^,ZFOcHfY51&\.f=CLSS4:8&8&7KFfB\(FJA&Z\FXTW7K/CI.
V7-ab,8dN?:6f7ZDYXRPfLCEfDI3=2c(QP4/(fPDG)#EY19)U7_99;&X/BJ=#:RT
E^[Me,.E_,/U5Y=10T28.IT[LZ.O]D4,ADA.V@]KeBC,;^2SRGVNH8OQ;7;6_P.H
JH+cb&e@O\5WIC?0R)fIDDEa\N7;I01aSCOYc+e)#VR@:[a<B)X?V^[MLDA2bJ^2
9\(EZ;T8OI.d=;0#?K4ODaF;L0=Z>;cU/:^=>)V8d]D).]2_?B/@TZ,W7<)CIFfJ
^XYA+3.Q07;R8Y(N7VY<X1-K3eZI;=fSVR8-+ETOFNaD-944/cbBBc-TCcM.C#[R
0e[b-dCJ.^I@./70>FKF\=PJU+X57g]2?9W8Y4#MF<SSDJC-O=&8/[\9d:,7FJD:
6N/U6RJ;f;f1UOEQP),(gY_^>0T0?8Z<T8B5.0N1gE0A?;7J]U4[&/L&c22W;[^+
2Y1B:<L\0-@+O/IMO64EP\&&UBYaE-/M8B-<\UUHY)U8F-X(81@NO=fO?,O=K4De
NVaN3A?ZJ;.[.@0<eSeO1Q0BF(N]1)bagS@M<bJD9Q+:M1L60FMA^9/V^SPdGQ(5
P/GDGP@E,#,fc[d(A03UAWPW02_4>dSE1,9(&(BYI(]7/FETYC9+5)HM7=ZL6A+G
D^e8eA]>b&]R9b>(Ife=f\CgY85HZeS]5KCJ,AKcAbMRcCa#QS>>NH^3]dY0@9B2
56\-aN;^E;:J(e?CQ[2,)G#F_aW77#BC7b_/.DEMXA&d9Y9-\=6a6Q1D^Q5eSTKf
+SK(-BE\UIcZ+K-H(TKY[940^X1aFJS9gOI\5N@de,P?VJgYR-,c&>(0Q?D9^@V>
d<TK3LTf/A831JT(b(&U0VM=Cg#],QS1;Y7Lc7b^7/:SF4^V1DOA(6_REbTPX5^g
d4gI@H(eX2@8gEHX=>eW06?N(O5W0WaR=g:\AF6-.SAcX85<GSDgH^6.a712d^@c
::5[JOMD_?f;eZZ6R_??4U6Q1a-fS8<57/M;^HUYL\)UIJe=+BAC#>\S9#H7MYNO
P&T4fJ/SEH<SMd\6_(2CV>U?QaUIHUV:Z]cCD:XM_Q9-NdCJF&+UaI)cbR<UC.BS
M+GIZTYc>?LG6D+b.]0B(U[6Dd](b/8J7Qgb<LC#]KO-L?LcaXcK8#Ha7-QQ]4&5
MNVNY(A_P_2+]Q412X[<PbeF?02>DKJ_5L\K0LeOdVOS-Zca6V3\34SSVN8BgZF@
G.=daP77b-4b@E/T^?VF34afaH:R_B?)e#(_Q:.aeD#I22,RO80-aWePSLUHMg^d
QI)K[U=Q23&_5&#[[-#OE78Da9PKb^ZZ4E[7);e^+fb9C,0PQVR\aMQMY6WVdX&C
862LHXQaBF/)E8;]=V;,9[DKd?+Q?B(8E]XLBfC?GPZL&.S[L/U\-7K(ae3H-S8^
4QO9f1VfBY35AB(]e&]aZfEV-N;X1L;):cA+2(,3^+M4L2cNg7e/2:H)&fG>_,MA
g=S^5-X]CB],F4K>;KW&Yg6[7bTWOQ1K(>ZX_B\7I^McVa/7DJQ#0aGdCWT2H@G,
BX;cLXV<J.4BY2DC>F.EPA;LX8>fDP]<]^I+C2?B^QSZP5;(fe/^7J>4?N=6\)2(
>5@N\g<L[>SfX3P1Z#KC>CVF-A8^[U,]&ZS+Q\U\W9@e5)<gP.N-8,4Xb-Y,[78\
?IT1;e-<WVWdW@@3@SecLDC2MVTQ31d.S2SE;2/(?8?307Lb_PVTT]Me?YN2OST(
KFMaJRSA-KKZ0XMR=MQK#HR25VBNUQG+X/[-IBMP.B9EJ3.&g-[)9TN1FV/03+c&
ZQZZ)Eb.FW89F(XA8_M^4)M^QUf1WR+6-/\L\X\1)g=UcdB-efV=Je[CO/eBcI:C
W6E8--&G5.N=[d;9MLJU<;ONbK?25N9S_fR7BF(@T^a>>1@210D(/CWONJX#IR+6
0E@Z2ZQ9A:.?RQ57BI@.,9R9YP84@AQAT4Yb-K/]])f[)D3TIbZ:^1Eg8&POefYc
,aB/+@\+)Y>T/0R;C)@aM@+,L7R<FQ-dCZ[BgK9RUDRAN[:01eX3fGJV5M\]@8D.
:<b9^c[SKa85H,3bQ):&7,9G]/[KUf6ebLFGG&bAL[=9egGPcKLeMXd?T>)UMS-5
GRJ3#A^G/&CSOP8\/EPg\[Z,=g5KWFH7G1/dB_B3E\ga(\=DaES[5]#5JYQM6J[6
fAgE]VV8^=2@\GNGgLN7<3-&ZD.0,R+-?L;5K,-Zb>cZ:6IS[C[/UB\<J5Z:\MHB
+47SVE834C9\^IG]]a9@6ECXfAK5FXCIJW-LL^XT5M?0D7U[#ED)Eb4MKRH)N#\2
.^DSdd)T3C3V5Sg/>Y<W&^aGW,4Q])==[>BGeA=\)_@Fe<)KHcD;8Ud^.:WbAI7[
+6cPcAV:#/#d^Te4/&b3)1H+Eece>DbUEgP_;2C<gg]@DTdA28fY5583AMb@.\G+
VD\P?Q9V_?9(XfD-Zg(dODTc6-V[71FD_\^W14.W>Had=AS8:[-79GFG2D1+g.>?
FW)M0:],+<2+EMY3Tf3NQc5S613)OVd+>Y4O;BW?HO8/X\]R)fP3KZQ&ffLY<RTD
d5NZQX,g6SgeZ^^(M,Y6gJef/g_.;YUbE3FRM.dAY8NcHRYgc)8PS0RF.#9VI54c
#?,1a03,0(TFX/E\ePM>bJ3_;7<eP#>g-K4(EX#KAUf,8F:1Gg0MM>6U+Vd^/\K(
5LRM<f6[](B^:6;KN=+>\:M-R@UGEVQ)W402VARRB#2\9UVMIB/0K=:&U-.M\8O[
V\&]W9g<EHT(3(8Wf2R&2PGVL;:FQJURK>K.dD(Z6_:K?-DO.YPKTAZeUP9BD-c[
V;&E4>FT2O)ad(^U9L]/HU-P9>b)HQ;gR]@VRR=b=<)]dOdWeaOIBW8&4Q]4YK[a
#91U=D(_FC^J[3Q.gS7b:&\QbB)T;RIX:T1:QH(5aN+?5+(R;L5(]ER/+b</a-+@
Q8AYKG2KN[Y@(.]MGZT63X;#Qg=X^g8c7\1O_68f,aZ6abL)]MFOHYQf&\fR1T[@
B-BMMFUdJ]g3>]RdbSAKB\3O5X;8AgDD\1;Y#T6N@QI8&H?/g11d-JHFfLHM:)5R
Z;eATUY+E2<d;XRKI4D<c)X_H0_>dD83=>#^/9C4]39O(XI#0bFdRF>Y3;UDDafT
AUa^N0M,3>UD:H7FAPOV.B=T9-0RA(/M&3KRY74f5cD5O:6R#bPWJ]2<<EB9Q]L;
QdSGL7.?QFeQCA\RM#A#&H5+_@]:V>/97Z[egPRbS<7NK/A;]OHe;fe[GXE,V?#S
[AP8MWB43WDX)>J.=/>&///g@BB0EdII\P)b9#EA=?WNf29N3L(+Wd>M>31:(;SL
Q/b^&R+[C)(=KH<7V?:9/8.<gZY;<O8L=<G.(J^J:+Q&QWM<C</c;)6^@Cb\8]FO
cb9KfB_8]aZ]]UI8+@7/1F(+_HQ[bTNG6Y[5S><^ZF-ND>1LH1Fg#&eGNZLT0.#L
7DXR@(&#\,+&dLJDMY[N(Y\YPgB@GHQKaC7)e]A#PON#[,ZTT/:_@2--@2MDc,CP
^c4Z>IERTFAcMbcH2HPTg/XB8<fM7?W7L09_38/9[C++JIcP@EUER@cW.5P/\(6]
AV]ZXH+L^6<-Ba,1+D(X^F0/0V=d@Y=@O(P(R[(:A2VW]H=Q>P1fJTDa1dW1Vb:T
^ZN>6.=5dEDFf41E:GLR-X_A\IECP?:NPN5K>.R#b@-NL(,M\/VDTDaR28(BdKS8
>P6WH,:+F?UC<UU&11V5G_1[(W0V28Q,-L[M@+(61eOK26Ab8<66>La;PeJHU#Pf
/J:&X)[4/9[bCD&7M_RG8K(g_B7)BaK=dJWI9]7X:JVAJ8(HH.#-Q=_[_3fZg-c7
AKVUTC=;I5_9P3+[?;d>>0?K[E@]/QN(SR,EgRCGc:=?1Je#E7F@V464,GCA1Ag9
Ab&g@0EH0S,19;5IC<FR),JLdX)CF)2;WSK24Tb(6](2c:\DP<agEUM(9WVN]UgK
BFMJ8W:e<K24&D[#,B##;1L3T3]P3.1@fZ7A5KY_G7caQ9XX[-Ya/]Ccb3>HgKC?
K1P5_H8=]G0G?GP^SH2:=9^L.-/DR;0&9cd-C<.<L.8<?e+K&<ZNRO/J@8TJfN)g
R^g/GPa<?0?dE?A0-&-25HQ@9)2=#@_-J9.Tg5\@7TG=56T5gQO&+;H3BMME2NRa
GPEO9OOJS[0B&P[VKb6N\_.?QX2<M@,)Z>]V1fadJ\5bBP)A#0gH=66C+27eN^bK
fM:74?2U(+#GK-d&(+;._<?NW;:1K(BZ#GCNL5XGUHG5E#N=0cJJfO0e43:T=,be
)_fC0J:(I;TA+cXa1WfCOeD:##\AZ5(d-#.HIe.3^56=+[V/95+C,<_R4DFD+J8[
5Q-#OU<H:bQ44/^>FU2gd8BW5>+=IM3L&LXD7cf8<N0C>&0>S?1N&YQO^Q-XW#X7
Se0_8Tc+_8A7O)T.U^[Z=-&&]H:[_S(O@.>L]aY_JIbfUA6Y\[>3+(G1FRBRTX-8
]LMY61b9\OcI.g)5FgRH>+RY#eL#UNA;QP6UYI7f;&cD(5[=#H;0PO5Q&32_PI,&
H+LGYa(;3d=J\3WIG,+05e?)04e-M>b(B,Xg8H\efH2Wf_QNG^UOMU3CJ2T,&Q>a
>Ag:_7gZ4<KaCI^8LCOF?OKcaO.E4B><A9QR4++>HCIcVU_S/=LT[IJDE#+>8U(1
=WMEN5ZGb#Q#??RAg.F.?.DcDIfL#-YK8;7bNP3/)QK9aXUT6QPH<]R<>YQLFK7C
aME0DW1:0fD(-,<3Ac3F>]IDMgRHc\KL\?/X8,0C:R9-RLe,/T)]X<YE8,e.@/.R
T/-;a++)F[dR6a=F1MeC75/]IVUf9P7Q.SBD9Xf_8W>L\V&/&MBL]:Rf5[0fa&C(
-QWI^#\9)Y0gSJOR6QO,Q7<7B:@Bc3V\57:/d4A2;4-2CZHQ0M_f4/;:bPOQ8)g_
S[P8^VGK>9YD-#E&gNQJZO_ARcE.b_aY-3bA\[I0RQc-P8#4ED,PC,Q=^R\8fJ(L
M,7&\Bf\PDZM7R]YIQ:b/EM1CdZC<^3,(DZ?=1VA9B;4A^e[1IRL4VD:[<ZcR:eW
Ac=J@b&7RZ(bgdDN,^6@fDA=9(gZVPIV@36@G+_-[0JJQ],4J&_-M>fU4I\(E(3[
.(ZN]0CJV4Fg[eB,3JE0:,1-4,5R#4V8eaZX_6QRc_+,H3[NMT=f8&L^\-g9cg]\
&(:\)\DHX=\fb6fYfVN,2Bb5U\b<3_YBQRZ6S7ZZE:L,^QD+N23CdVP+.8eVCfBc
?QO6FYRG@PKMC[^e&a=Q>10PW#=[Y500V(geS2.1.^]PW?,,1XW4#Y)\S]8L5)J3
5F)H0KNPM?P8dS+8;N7g8R@SWPUGD384M8f#=c(=NF4c,9#R[GUW<d2RVC(FN8+K
_\6]SH^P?VCWLCT7];_)SDQ_\F/,f#N^@ge.7\Y74M0X&UcAXX;]9-Xd+Z1JeR3_
6P@cSYDED99=JGRJD;(^bDP@=,BOI)W;]9D_1M-&#(?a31WM&Y3P\-Ea?;XcA:C/
YSdJUL=B?HY4]6O61;C:E=,3TJ+eP=REG8gcg[?\]ULCR<_>P):bV@cO>[VB2Qd.
KUW_<CcI_J)-2JBKU9906\:@]VD>.;d:dF@VE(RF@6G5=IXd/?eF1Y[JeYOWY-<;
U/B)=g8X9I2_RCfZL>8/Bb33Qe7cNL9f.5T1f_#9845\\YGQ@0^e;MHYBBT@2e0<
XIb/1,fa1@V?8YLg[,I6c6(FFDO(<E++ZV3;]2B:ag\\X/#B(X/SG3f)FfATeX.,
JZ=d-SR6M9I\99Ff6,a[I8+RN;^GNLFA:cI60XcC8;64_3UD)@+\)L:dPBc5QFIW
GHO=[8#f^KU,/[#eaG^BPMF[Y.Zb6[#0?<^#S\W5VAG(2RdO^IT,)TXcLP][^_+]
Y70450+9ZQ^\JLfZ&1MbaP1+Q2ce(_(/A[NBN5/],074a>B=bV2c3)5O4_D^-32A
e96_TUbU8C#H&8a876]XZ7ff:201_3H,&+@C,[<UG5D>3G]PY:6Ta&Q6(0GL5-0P
HT@;R@/V/RdL4ZED6=Pg_:EM)2;-U1FANcR8bL8G<:IJfI\,,(LMDQD4G.cO.^DI
GRd--X>cTef5FDbQF(>UFaVLZZ-cO[C]+L=g<UQO?:2FRJaOC2@+AX;c3]_TC7^X
Y)YWYKg)Z]\)[C@/C:L\:K6Pb85ad#,N:,-KV:54fY96II8V)3\(4O^9/f1:S=))
1DKG=WBX)@Q\(9KfT)6f4RNaXeR.IF]Od_&<fd:#=Q05dFN6VUgDG7:3\=3OJTOc
PecG.C5.RW)1Z+4E130Yf_J>@>,c&_>[?=^+HU>cM?ZZLU@[,3(H^Wd323E)7)83
[>M1Z^gXM68V+I#JS]dCCd:GeG?8<>fBBfWQ?=aXBL>KR=)AKgeHe)FWPI.:_VT9
cHF:XXI=U5H_<>ANY:X9&;_;Y-HSS0H6B#D2[ZV:^g@SF6,g6dBBHcF.#^9J+WH,
2de^22NU@Nfc<a=VRT-B)#F&EWa]c0G(Z0aT01=JfV&\C>O[CBDTSX,72aBN.KEg
f4QUEVYZ5BA>He[RP./3-4XFZ>NHO8M5R4WYOS,(YRQ@+KG/Qdf3YUH;A@e/(>)a
[W2K?^g\#QPdG:?22KC(5?G]>PBDCA?-INY[YL<g9O2:gPJJ8[=gdHQb3<J5L9Ke
;g8YPS+BUYX_]V&/e@U]&KH3,TFZ;g)@9L;AH/<3XY&V.&SbTa;=S7E;>bd;MZ#R
WEA;077PX:/U1)9I]E1VfNT00HQ017>0M_[Ra1/<]:D,;-A03UQSO7:0.g5D>&dS
HH+FAO<J@=:7.]R1L325V]U;840S[:<D[NWDX1??P7fFS^QAeB_+++MY:0&I/&);
WZYG7U7;[ZQ@I8?PJ>2B+/Z\_(2KfJ^)4C;1^>M0c=gRSG]&1W;8-L;4<W[1&3AX
U,;_fXDOf.<F_:JKGYAQS05U8TJ4L88L]^-Jce>(a,^<6-IGeW;,B=([e\CEEY<R
eZ437@a4c1.MCT/IfD4NCJ5H?R&e3dFKK(?@2/Ka.@_^,GWfc34,:E6#c&@,B94X
S7;QOaB1/>CHb2<g:P8]T(G&IFA1UKBgA/WXZE?ACf,_PXP/HY+K#V1I5#[Na00a
7-X&-8b425T13f]-E-bXA/RWW[#[:O0CFX&MFLDS\+,UA9S;U#]-6V3\XU@/7HY(
b\cH2OD/O>J)[N=>\7__\c+g?KF]W(SE5:^1SPJT)&96#_@?gbS:)^4^C48/<<_T
3#&ag^^Xg_FCJR4RZ;\>H2cf]9JIB./+e,g-]Q78HK;2DU^#ePW,PM&1g/eA<R:;
5EUVgQ\F>0QJZ/SV/4d#+3XM,Ua=B(W6H#Afa;&()8W0e+Y_T&dAZ8/:dMFGe(:&
ROVJ^#>RJQ::c\K<:YP-+LXa#JKgGTKWWd/gNXTeQ,ag59WXeaPZ<b/WUBPOSE=<
T&V0dH0@3Q&_X_SQ0S6AAH7D)9-,C.:b/M02TH?HCWP8.BD^6=<=00=OX9H0^B]Y
?&\JI<3=H(cMW==M]G8+<Mc9<K:8dE[\3_O[:Q>2T>VZ^g7/aK7c_a3M0(3J-W9O
7f,<EXR3@\LP<O2F_;Z(TeHGB6_B54&[^?[@DF#LVc:/0NIWU7Q;Q6R>T?fUW9U8
#(XT:LB_M<5M&7DL2[NGCP9fH3NS9LN^NccR_RI]DX[;4aVP:,]aN9WTYNV)8YD.
+81d>&3aBQSWMTR42Eea;\8f&BOY02KG1Y051aAIS6[S\\HYQ:FNbC+0<WU41eJG
:Bgb\aT\[^RWL@NQ-NM0061aT:].?0EWAP1&#cPK/3_OB#aeG;EHLZ_953/5F4Bc
R-K)TSIN<UL80Q0T(9R6P[-_,@gA2K/W76Z9PEDZ?_W]P@+;#)@?5F;.+M?4[4U?
0ad4<=\]>[_E5cG-=/e=c,Yb_HFSc#]I4041+D91ebfW>Z;Z<)^/>=;Pe[(/[cd:
.-2+;(@AB?CW9LB1[P3_fY1\.MOVY)>EU9CCAfI5S&X5M/+B:c:F71)bNFOGA^OY
[G4.3RE3_g;8YTJ>(a71-0<JNe8G[<(gXWA]cAW=A)_E2H<M4EE;P3>DZ+5;dGZ;
Q?[cOWa^)cQI&._,3(>_49EP>2O_2U)\_QJ4g+E@;(5_8>=+6(?+8ESB3CSG9VW4
:W<)U;>:]TQTfGdCeE,>9I4>IZI9(g_]a+M;5T&MXe@(]TO-?6<@/O3GD?_P3<4S
@)[R_QP)QV00(I,Y(4],9fB?X<_>T3)A+b1@)]PIJeE,F9fC9G-c.c8K<4f5>M<f
@R<5Y;:B_J3-?Ec7K825gE;,;822(BE:&ZL;IXB]?JdV]a\F2EVN\1gVEU]6GLK8
G=I<Z)RBBd;a???0NQ_L\OTFN^ZNS2Z+MU+3^KX;H,dA>E:[)II5bfVRHe,_Lf9.
D^P0fWPJcS=gUd&<aaP.CVOg40.L;<E.eB/1\=>VUZ&.A^7GT)Dc)0J=\WW1He0[
-)0[ec03KAURE_42;b+;1)g<VRKIJ642]=AF.2EVP.Y4GP-#E^3R/_^C1Te-79M>
^&:=(0Q].9ZU^=Jc^Q0eB3V.BI=B-E;eg3^PR+TGF>)gZH:Uc[(19MG/NK8FRO^/
;;;:Q^e:LHH0ES,2#^d)(.BdMI4f?<4)OY\SaJ:XI\SCA7Z.4R3OFcdUS.#L5Y5.
4NcQO__OM2RM:]70W](7W)I(I9A.P5>NJK3?YBBGaCR-W?2SXf/XU0_:\GX=cU4M
fcQ)Z[D;b4>Xa+J?K8g@VA-=b@NVRSQK\=^K74&6MS(+\MCN,[SG/>>AL]\RO0.,
)QWG/aG,^>SW-XL8TZ6-J.Q3TQ-IEX:9@Yc3XQO[=RCOA#<_]^Abc<W(GFIJCe5T
Tbcc?U7?[NdFX<ea9>d5G6N@C@)d#JHE01+6#D72<R&D[W]>63X0UfSbU_B:aXWb
W;C[\WZ6/68)0/PHBa,M9IPD?<8L/5HR(DMR1>LY_6<>F\US<UJB^[]ZK^BD=@BU
_.S-H>?-ZD+53M_6_P+O@KCD2=)]]5Q#:;+/N=]P4F,M&Y..SA2[3fd;?M43OW&^
=BUT:6:Y[;Ed.aZeOW-&98WdYRY+G0AL5eD4@.B57c=P5SX<V1AC4a^e:?^_[[;+
<@A^LgJI?3EbMC=QR:6OVL<(@AUT7,X?,Z0]\S&;]d_L<G90BYdbRC;0P.3:#K+Z
IeC[<BN,O/VW\10[cDSU@B(EM:>a@QPP&:J+Q-aVP3BO.;E9@@GXA#6/2b32DRb)
.]]I&_M;^=Y=F]c;9adP.MIAPI4M_)TQ5c0K6HB+LId.CV[(/Q3bARLCAANU@B5Y
e5G&7O8g:/SG>ZV.D1;^.U<KST.3J_/_a>&)e@Y;)a6D:P)Vb2=F>[.(f6_bJd8)
G38g3QP>N,DUa7+fR5BU,I?9K7/0FR^=FOFYU.4/B31OS^RJ,]g,@F90R9EPL]fE
C\XB)_dAK2P;BB3dc:._NP)ZdC[#SF[[56PQHMBYVcGTOdNM1D<R:AG)9O/M2I;R
IWHU^@;K=JA?cU#WKR(AdFHP7^?AI&D\5]A5:/G(5cX4JI\Gd79](0?QcHU\I_Y6
0V>67VY^FL3ZH,2_8\cN8Ab:^C;8A=S(??S&;Q70>EC8CUVI8dN.D.-d3D.8)\@B
e#MD<T36Q[C;ZHb(H7L7Z=e_T:+IaM,I(G&1;JIY&8<B8^#L&H:+>N;6K+ZWeg6c
RgZ9LOR)eX,SJDg]ISZE7&3E<QGF+)<7@(C5KgG_G/EU.Ug:\ZK_X^3@5Ndd7FTF
-+DDd)##2618c@Z/eU8-(9BK\BPNLc,.H\L(7HS=WB6\--\779LUHGQZ>NIXAA5Y
Tc8V7RKEEc+,;a[S1K)+<J-?L,e]]Cf<5TgK\?OLM5_@HJWEg2ID1QZWH@YI].Y]
@aZA=0<?#2:HcDTVMM??PJPG^0^c/;JOdX>bOR;_/&><7X0[]00,N-6TEbKVC:9P
ZdYga0WZ_-0)f;H9bRF2B#Se0W=5M-5W7TC;0N^[:Y3]->LE<7N.e<SIYDe;9Y7R
C^-VE3fPC]PP,(GG3P,bb^+#UEYc+LGW25;/2H)6W&ZM:,/C77_2P#2OL/D\7_bA
FE.Zd4D/.9;A&W:X6L#T^T^f2(,H1,O6e9),4+D8DYCI(8HUV_/1JMMU)F#3SG0F
e-d?0F(+47@8&CHG0]ZaE5/C7B-M.ZI&VP&(>U>Q4FP0J4,dRC,<9#fYO6-]O.LX
HOVBM-Z+,]bLM9?7<4VPb@H/M.4M8/c:1:6/=3RJX\aWQ<g(EVW<#;)^4YVTI=(,
A.aAVS3KQeKd06GA?RCa^]@0gYY\YF,BCAGIX8d[,DQBCS#^MT)W()Zg=+(@X3.d
E,+4U_ZJe<\-VJ>A<?IV(:d1gWEU;.?+bXFC1MVTX.#1MI<:B6\;6+XNfZe?b2&+
GH4=.g77?C?:<YNaP==:-(\^&55-NI3]OKJ4WDdc<g.+gA+2X:CA^fY;DPaXM=[Z
2^UC9UW0-g-41ZX40JZ6IHH3d=+X/5\2J.&#K^E39G\#.?:(I99R<@ZdVdPb#2K\
+3>,:=d8B8[dT5WVb)QDTDF8<YI,:fB2T]d6R+UJ/H[C6^,3_Q[2aUc,(#ecCR;Q
Wf&#>5N3fQD)_F[A4\2;SIX+72(K/f9.VBV]7QW0Y?\]6#8A:0R+YKP:X<cXHG2(
W1VN7RVTK2f+TX^K0e)fI@3@M[/+VMF=DX>8aZK??R\&VB&QPH_QW6\V5NbISF)4
7]-)+J#XK]0(HTA&X>Oc:,:O)c5&;-(=Vca7_c/Yd>?d]W/d+78BU(-\9;X[JZac
QTfKKF_MO&(WY?J.I817B<aT0Y6^1=E.+_?Q(&F^_W9+&g.9YJHI0S4D5b\/_Pd6
VUe1B@Z>c[.:&?D7NWde_D_LA<fc8;)F\D7R?/9@@d>e<UbWGQVK0G3RR=KBAGN2
;=aceA)Z:@WG#/7EU=PAY^RgA/0,#EG_Z[H4>Y:#?P0gCGT8XeUDb3_SHF.g3JWI
50b&TUb-.1@,C(X:W_fV(@29C0@I3J],)=c)IH1D74\b^.Nf<e]-[A(.ZQ&g;N3>
5C)WfEU;^Bb=eQ[)_@O>H8PNaSM(Fgf9LY;3b@=W5R@1FT,I4>8Z6/dF-BbOcY0H
8&\R]\OXYfA8MF6>H4_D-4^\f:OU=9/9586]KI>Uac&fVcWFWUB.,>.g(cc@C2HD
I0a52ND5ZJG)F4N(JZ&5XRbZ54=eWN>QOEP/=:8JB=cJM773Pe[Qg]0)>g23/e,+
YM97GP&H.X+(Z@J.\;Q(-E32e60W?2aEPAE8X\bHVS=VdOfR2(9#>_N<LV)M983^
6C+#NFP_IR,E+d]+Z0(BD2TA;KLADgTPX@45YJNa3E;IN4;a&UI+NAVFVZ)>AS67
Qb;KT8^IHa.P5T?ddTdCXC4]D5b]7f^EfF?N]1N<O81IOR/?9[=5UN.IB&dS&FN=
.g#KJ4+F_gc4J=F,1NGPV,7]ND(gFK;eYIC8(0Kf)I1=8ea-GN.I^ZJED?+0A#;&
)^[3G,WfCZ_]0f[G^;Wb)3P).Z(PK-?=PB]4DDZ_)D)bIC&PTZe:a^C4bXbCWd^3
:CM+XcKb8XVPWW+LZI@?<3YF/#5PTY<98,dD29-c-NAB/GHFI(SUeMO+F7g@O&)6
)ZP^;GgLF7#^X89(J9fHHE25dIVQ.WB7WN)QNPQ0_16<Y+7OcEg^>7<</:3L3WIb
GW-Y3S38Q^8CM+)P1GdT7,,bc8aRVLIGEYVQfKQGS2UO.)O,I,)eUME9+79H21)^
OVFR7RS=Ia6CDb\H<7I&/f/;;@DA1L:^Y,UGe1[->KAF&WgMU>Q]R9Pd@5,AV-<Z
C4E9H7:a#,:(KV^.cZbgAUAH=F4A>]PG_HQ9X^_O1AVb+5#Rf/S8RUSaDfMU7geG
WY&Bc.85L/U8JG/-5F4[ER,a1[;8D0+W>0;D)^N]2G<5^VY1CP(1XO9D>7QJV]N[
;5Yc6]Q;Y4Ib-ZYIA,MSd<a?EL)VUI_KFCAc>b(N&V1&&W#cQMC9S5&(TT#HDP8@
O7cW85RF,O,]Cf_Z#T?2/dKYFT64@4R\&<+<9^^126>b?TgBFSaUdZ;Y-PIDLDKC
.;Q?]9M3->[FJ)44cR>FB_UI>EY,9NO:/N0N3942[22IVYB0&1HBS9R.5QaJ>QfL
WLJIb+fAIH9A08;TA0aF&J3:-Z17CXbb030Ebf(G&;PD]D_=:B&]&8=BJ=JYS_4#
_&(-f-Y<f&c<-5&-[)N3.He36g>1eJSV5QZS\_0C0e#BJFagUa],RX9TGA6UdX;1
J>.FBJc3]@(fX@DaT7@dN_IYd]6ED&,OTWRbE-e-JL7D9-L=8KUCYGbH#1OQU=T5
G&DU>=S,?\=fc.7d1d.\O/]C185?E_Vcb]bMBdC-0W>OeNTJ47P;RQeL?EI9F5QB
[)4O[Bab\(K^9C:EK>=Ke<Y\8-5@SL;-WCf<EZE0GbHNI8SF/:#;./Pb;?AW)W@.
&G+(5ORBHXT3bI5egXCTLW;A;=faXNZT^D^]NR\#4a5.>a/K4)gBRR-BO&8FQ[8e
_/-@&J+A<^]>U?J89N:e7->+UA^NH\AA^SC3P?T;MZ&SaC,R>]EF--gSYY.<T#.A
ZBR[E8;P,9,YM@F2^N&^B.)K>W&G>P?d_ePd]3^F6]Gb>-S-D4.9Z1g7g[];JWJb
(>70F7YbMWH);L_7Z\DT?<.?FEB@-8S?PCP[aW.P6/S_c#8_edB04b&a_VUQI_1S
04AUNA>C.R@&0TN1+a6-B@7T.)+/O;ET1]GN=]R:8aAVR?.PH6?1VLGdW3b4LTaL
XSb)12K4@GTF@,AC\1B/eJ<R5_DWBS<E2&,9MIECZ^O>A<H_66N+E>A6EC/\FK#[
AQcY4?O6SdZYK?@Ng>^Vd-OU7Y4/+P+LFV^()0^H8B^YLAXeKG_b#/83]YZVaH,A
JMb4QTK7/JcH6P&\\&6H07:-\eW=MF/^](fK-+C/5>eP<VY<X\6?&5;48\LO>:SN
g_KP@CX6J<3I^D1DJ<HGRM/G,^7dU]N)I_9UVLDV,4=;4gNM[)^STGKE>d8;OE0N
,P4SOY\gENfb)0g;e-IYQNR9gc7YAWZ[)1.Q/f(_?aAKZ9\-SBCO^_Y00W=eY-GA
;8[fc0<NV2,-d7ON_[df/?fC;OE1V8-YI>Y96,@d0YU@)0K=0G_ggD[Nb46>?A#:
aIWFgFZ-,\6dIPd]gDPQ7MC1,WSe=@W?LP(@\CT[AK3IIY7d?c+7f30<Jb\99eY&
c.gK\VLa1R6)0PWY688JYK@:aR1VF++-7SSBF9SRJ5L^\Wb_e@)IQ_<1U]31.0@B
;/CP8S,;,N.JSD])0CTa7?dK[__H6>&NS1M)bWI^C^LO1P-+X3\1TZ3d8F^:[)4E
Y@>GcJA_=cO.FJBD@,fAb\8:AMM-7>YgV\KgN)AXQ>dD+#6PWbgD]4+W=,66B-OJ
#<5WLL<EeK0J?<F5WJ@c;XUJH?__cL8##HTWX25ScXIP+-U6]?&.W.U&W0WV>KdB
E^5Z4RJ]+OB?MM=]^c3=fNT.8VW0NW]-TA96LR&68K7\9QA&X4PK/cCE08/UZ(&C
.a60:GK=0J).J&c<7A)7>Md\X61T,CC^G^_M&dd>?^FO5)XPO0Q.OHG[(/>DET?9
SB.(B]>I>HQQ=ed8I#?F\]\\D0S6dOY?4e#MW:/D48-(22C8+aV_(Fc;gNHA-^<^
,ZL9]f>+M&e(3LbfR>d2DFEbV7K;+>+__.3aU>6\e@=f3M75K572Q\(,F<SYRL&>
gA.If/<OQ+2-JM+VHc-[8Sf2@?D>5JTEXWZGCL9L>J0]Y;YQ:<=^/SG<S.\1&_Bf
=3K]c#Y@K^_\B_4R655b^NF&Qc^8-)^,CcXggS&HbU\K?JDHJ:c/@KdW5LZ<N\(;
+=634K(R^>MP[Y;)6a>Z^G5Z<b4c&fL]<BeEVT;=^:8_SWL&2B19Y3\8_/G@V4V?
=>gZX,0?H#,NM7X_&WXD,/Vf&^\,ED5H7XZ+\XRVE)LX0)Q(ZSWdXC#C;8=Z08dY
0?FZ+1F1-+.ZNEU;H=J\V_,?ZKGg1.a\73aaEI]_8dZ;]I6/<PV=(gO,#1ME-G5=
SHbJfUE9HZ/f=P+9XHHa2:-6L=]E=9DRbXVGB9TYH,7?8?g[bCMJD)g+[D3<]X[e
OVb@8FR)Z=?T,1e/b]84&_MWWH(USD32Tf9H7TJ31)N&fV#-2(5A_-U,AU,98V<=
Sc1f>N=FBdc[,Pb,WG@U:a\C+1aQWXS4e\aMAAF<#V8]2YbagQ<0CW,_?/=A2U_g
S0dC+_[Rf.g?W[4X[)U23-&OfN:;O,BQ^QQO:b=#8d5<L<.)eE<>a9>Za)YLFUPK
J=?TH<;)9PF?[<.2X_5O5SR(=1O5Hc7F^6G&)d0=.L);061PY1FMU,Y+a^_fCS_R
)QB^_aF9c4IR2U)a0c+>7-6W\K[O(O5PO,cSc^QF[_S(AO-N/AQ]&WFP+[O;Pf7.
SY/?9Z1.8-KV&V?,P#3&V1)W-)[3EBG^RFL6geZDYCec@V5fAHQLTW\6WVI3NF]A
CZ&FJ2.;5Z)EG#?S\]=/+0>UHT-#E@>+WAIK3YHgR?&T0K74&10Y8+69D=QPTRLI
2/G8OTDAYU23TZKcKX7.MegGYDBTR8?.ISEY;5BVF-AOYPDae)=Y9b_Gf,_SRL/K
@X6BTU+D&5WK9a(D#[0=E(gYO[:N,@NXd?\>8PDWTC]_DN+\[c1YV000bCW:6Y&&
#91=;6bM7.3WRc]8P;MA)).-?M1[@#aF:FXdG4?NK6+EPG#UJ)YK1-WGF>_YVbWJ
?7X-/e\WQ;0-[a>0T;\E5_/5bU=K:\7Cd8/GdJ=PC;e9;A0>H-V\W72CXfIK/MG_
3(M:UIAa+<56J<Va\3b+02LXPH<<?>e.SPI0BDJQJY[,&MMI##XeV=,IdIbAXYET
.9J4M<6<E#BVf6[Ac>##5<?FONP6g-@U]g=-NIO=9F(H-@S7&=LTcB=,V6U/6bHR
Ef2eGdGMaaF#>DX#[ILRYd3X=D2W+Ug+LQFY-F;;_?fKe2&OHD&PST14f4C>OP=X
e0W+0@1dJ_D;9<aXIESPIf;e;N7N]_EI9BCY@@\IFU\^MM(=?3QI>=Ue&3\M>HD=
Y3NDJTZ45^1UR7@L^<=aIAYU,0<f=b1EM+^;^--VA1BBZ?3H@HW#J,:gAF&SSbDJ
HTb31g&dM\#[:\:L)7VFX0Y<RMBWd#AG+VGBVAI2dY)-P.g-@&#E03f[GUSTLfDI
/A[4Fb2[4fJ>0-A9M@BObVBV<4_/,gHL_+e7:7CTH/9(3[D#,BE+f.eED]L@9A,]
0=07JgMYA>6J^>9<ZZPHYS13^A8dQR6/A9OP&P+5<=GX>+3(<?PQM?1f_4=Tf=^/
>7\_7Jgd9U-3?[8B7C,-K5ZZ,XaPHW6Z6+HHRO==AAF:BB:GIZJLH<.bJJZaXBXH
H4PaI4KGG3ACfO3IdI_/7=-\>cL.I1Y?__FLZd40cdS6UR,1)&?fV/5aP._DMT.e
.LFgXYOEXDeAE-\8ZY+I)E++LaO&Q-T6;?=c)A-<5XeMMV2-R[,[VS6S<.4Q,.c.
CNIC+7[+6SA]#8WgK/b>C#QRWfN(<(f<c1)EPX#Gf9:W.0gW)P2Y\T;1=HCQLIC6
Y[bRMD0JO6V04c)?20IESD;O_9]?Mf1O#K0GG&0:YRT\K?8caKY[/ZN/bM:Fb^Kd
XMRST1X[b0CId\3BVS-Y-c=MX)B08Z.Jf:#M67e.TMM3f9HZc?BK].F\6RY\I-a+
4W=6VBLI6]V_F9+GQ@d.A;gVB0K,b,CN=X8R#Ud:a2d:cTQdf_W+.E8H3_X,T&d7
KY<7KCVd;2>[g)MSONDB/f&5VMC,K/-X/9],08M^?(V#;;-b6?>(Bgg2Z8&NZ<)S
M?b?5UH(6D\EW-N53[[)K98Y=<4[^3#Cb+_W;@TPZKXO3_YaB.aY^JFO0C(Dg(d^
GPbb;?9&HI\JGX]6RQ=Yd6XT>NY;JLU(D35ORS5PZOPGTHB-H/AH9M]BF?a@WIAC
CEaP\6(K>5&S)_>G#b1=@KcR,.;04(gc@^^69)4=]d;_a?VQ5b\fET&gBR>DdA9&
9X/NL8L4^82]fV4^d[WB>Vf#VWGZK8ZVH2bGaIN-_0N./,5K;VgTI&R20UU:7YQO
a7@R#/?8b>.53H<E@-7Ia7XM@#I[\V,Z&216LF+SDT&08H12I?)Q+<F/\7]U+7.3
=.(4eeCIL4@B)592)>;<dJ@.a]8W-O#Tf.CZ4]@T4Z+YZg7)1.PAa@b;e([=>5@(
1^d@Q(:<.RHWGME+a4g6gITd].V_Mc>3#5eTL>Q[2:SJ89:8/^)Ka<=?@T^NO/+Z
fVUA@-QaMfQ+1=MPML4ZO1f,WbF@c>8fEFG:.V)eH)Q:YUH2]RN74>_g55)d9JQH
?6+S<2a^]PfADKT2J5TcYQ67^KDg3GfL-\;:Y3,;8fIBfe.=Y&>-P7]fUK-#(SgP
JJRPWQ5Ha]1/#-3.@TH1Z>.>-OUa:8Z#6@82D.B@.\<J5[(c1=SPH7OC__/gKd[1
K0e:T78:+=e^cL>VAcW(8OVQZXBZ2^;5)ZOS9.BH7eP)&5CVdE3F&cNQ;&8&)T,Z
JI4\b@&-0fAc/8b8^/P@L@Xe8Zgb#BY:P]^K,6M+^.TUZ@c4HD@a?cN3GZP]L=D/
S@5G9M#28JG>0:1AcLGJ59LYF[CERD--<T)QQ0e-N89TUSO4F@0:Z_O7&7]+.a#3
-g&&e?7]2X9?_7RLaBaB&QIVOec/6Z1WS.RXdXG1=(d6BP@EF^>C#_O]P7dTg=-P
1NY@_0[LO/&fV1B7MD9-@<g^+H1M^<Z,L_BP9?0)]Ya0&-JS[A9C=J4.<HBQa&Zf
cc_8>1.O1>U<C3b8dfD]WE<@e,+g252\+?5DdKO+9,U@Na(]REIN@(SRU8_C@4fb
3Z8-#_QI_N.K,b^M;)?ddUP8)WDM(,3;.2S2fQ+S.+9.e)7bJEEVHS)9[#b5@0U8
>)KA+9d)?e]<a?[^+INbaXI4#6Af1\+EdDW:;6cUV2d,LWG4OKdTV5]ODOQLG>.g
1YGDZ\/SXQU6>=/PHE6M.]QBE.4R(c+Q,63<A/11K2;27#A;8c3@SOA1A.cPXG3Z
&BHFe7?V,aTSWdX>I1F<G\FV=\[5;SV)=>4\JL5F+7#WNU?Z2(cD#Z]]KFYDgCN&
2UFHL[g9<5a(c&_Z@Q(TEbC@GN4G;AX5ZPC0&IPEFgES/+)@X25J2N(WD^WUM5[L
6d=VgL&6OTW^]e=^7E6,N#\,6PfHF<a\X14DbYKQDUB?9-R30bH)>&CBUBGZG]XV
:+-VHE9HA]&50?2?.<FX;Z2<YQ:[)+&Cd2LAgPI>(A^9Xdf)>R.T6T3aS97=J_Q4
=6--PHL7&)LVL11DM3BE0J_\RNX<SCdCNOYI),XCg81_Z_1g&<_<IV0CHD?KcO;S
8KQ(-P:/dUcOKQAZ>WdKG^Vd@R53RB<WPR0KY>ER:agO?DcLH3ZUNA<JY?:L&D9a
<4_EC9I/[dW=dJI@NZ^fN48ICg3[E1-MEGLbP^PI+cU#RQGCG5N>fc#(1HJgI-C?
86VN5X4N2fa^(5-gKY;&WWQJC285B?N_\fF]F1^/:/=?_SA,927<Z[e?G[gL;ZKV
+0&G8d0QKe+c?Vc=JeIQNCgdROe##:MWdMOC?<O1@QGZ7&ZW(VO,OOO_/I@-8XBW
FPbTG+QY;-@Z/9=g<]5F8D:(BH6f(eCW<1KA2LX:dSa_]\aaB3WOcHFP;1YHI=+-
79(^G1HF8WeF6<ZFV&SE<>V&E1>P(?16Y5:gWGU,L(J(SNa(P)@fdWg5/G\gMe>A
IMP.&W>Z1BSZBTFPUU#_QeHJI1](@OaBOdOM1=(Z/YJWYbJYQ)UPUGG2?b_LLF6<
U[bbfMLPd&ZE_Ve[@+2\571V;V]5K)\UC)#T6=ABdHfdNIG:VGLgW,0Zd4=eKW0C
T)@KW)CA?J5L@]@(08:/RT#Uba.S.dTO8NgCd>2UeBe(23GH<KW1Me]_8B9J\W_^
0OOZXIR0L@J7H=J[Z+>7d)Yd]UM-]/gRM(OYN_5K1JWPG+f]R?=cNACB#LCM-N+E
?4>2I8c6D^g).&EJa-@=7;ab)b7UYO+GO4W&MbY5;d;\->02aX1UG4B4B17#FBF-
)I2FJ5L2O@+=E>79(Z39B:EA]=)9?P[1_[;Sba2LXD?H+GL,FT#GR@d@78OZ(\O4
7T9-OZeG:YQaQ@;Y7VKD=HFH4R(TVbGT8()+a&^>6,,G&;1GT;,37Ec>1fJ5]79C
1SOe-QG:1CHMe1&He&aG;.FNY[.9GL^/.)6/?gDO-WN##H-]5KbMHGNQ6?>E#<.S
?9O2EeZQ5;M^:)YR(0O_7=K:=76M](DGV2J7&[X3@4G<_+?7^97<_&OR9bFeL?8&
HfF646ACK#2g)>8P7PZ-Q96VJNNd-9Ga/T;M=Facf:.^WOTQS:c?H>J+6+dJ]I0F
3/#R7\)NJc#&POFa08LI7FB><4f[d.VY[S5M]7:I5-G8W(=I[=6dF+JUJI>U2IeV
#XRM1IgPG>[&(-@N.RCQ]LV+NJFO^C)5W_8e^S[#]dg/RP=YB.0MM2#(/4H^L\<(
2G4g?5OfYF[3,:TG7Bd1.D\?K-T9LBVWd\g_Gg+I])3Q1AM/0DJfL?2CMf#ReQJ#
H+KTWH\DM3d7Af.-&2Gge&_L8>T?^^1RQCJ).^aP7O]K8?fHE(W:;R9I>b.QU30>
@YY(He>13/P5(D#6:HRD(ETgaM7]>Qbcf<-dN#ccG.32WdS.>GLJW]gV#2I(5g6V
0,^F@L)F9-_OCaHS@]1>4ecRdAH1[C+<ReMN23/\;E,4g0c4<eI2YW))XFDQDCC3
.ODX-eO:?HbO5]=cT\&A36Q4g0VPN2HCE3^,9P8)C&X[W,W6[KB^B3_^-=H7?CIO
AB8^a_M14eI,E<A=YcFb3S1]YLHUe(fED\\O@-#b>5a?d/@36&9<P7N@TI31KA2[
Qf_7\K5g1R/=@ZPfV&J-1RP>.@@caMb#UOXT[,Z;@B?3c^3]b[45:7RT/+5/>?8X
Q1]3UP[dD==A<.=NfDB7C81dL2Wcd4=O]M/Z&\dKFZeE])/BEO5XeW)f]D[^R>e@
KO,[BBZ55W\86XVQe>&VPaQ82,_/FJ5[9@O)MY.-=5/A]Dc8\L)U:4Ta(>DP>;_-
/C,T.UU7(:U#X:)g3QZ_eJF1_^F_NN\U/>VZ,#&9eEXReW4TbVde99:@9&@;1MdX
2W@M7#>,:^[C3BDR+X0E6^JJ63N=2RR+JRW1E/A:CMKVbRK>&IW@1F7/)E&?8b+B
c+DB^6Q1)DY2;+2X4AN<d/<UMAA987RQI-8Q,f/8.1N9@c0L/^Lf\4VSHSI[f5UL
IUTe5MP>bLN4TG(6.^90-0<<QS_T0WW].^LHd/SY.K\E(ITG&FZdM4FfDD;^+JA>
A,:R^5R,8a_Q/B7-KdS-JdV[GAT(\@_F&g978g#I7.dQQ9+YbAD;2(L1OJ1OGO#X
\f4S&&722FF)fe5A<R;fIWSN[E4TWXHb54+&RWN7VY.-bPe<D>)fACbR8V>:+5JF
f2];USfaU9.JX.e??C..;>0IYLQfWeeQOIcL^=2Za<2^g9[Rf-=cc:Ef@60KYS/\
FSTAK[H]YJE]A,XXT4AOQ(,(B\ZVH,2(820L&YY:,<cS5Y<@:@JBB54fgRf4RFf@
c@7CFM#;;1:^X..#\B+VRO#]E7RYG2U&T@+;bNG^93Wg@#T;a;HYNd]CF&-(PQU2
6GL:XTR/K#DV:&C#DV]X1H;TTS.JUeHF3C/fMEXGU)Y.EQB.Ja/RbBT:7L=d#23f
\91\D#N=S>Vgc:F#=>b&(I;4fA_^b5NdCa9F7&G[eS+(88U)1\P3gY1OF[YK5]_(
AF5OA33Wbd@[edJUJge_fZMWLZd6:L\6T=0/A(W=68(1_M]ObBH&,/eDQE^a2\+<
aRW^MR<N-MA:;53PYP:Z,K-IKI8W_2CFdKH8UONG?MB)FY3.K=<K+@[PdH>MgBS<
NDCbVY]<IA_DH[S=^8-fFdOe.]f:.Z\ESE)[ZKQ:J]3Zd5XK^[)K=0AGCYfVJP7J
7PEOOQ+0LcPRDIY:a&?J&aU_WeDY^<1W<==?CXD_WC.d6YX&@;H--Tg)MZc8g^M.
0UDK.:XL7295K7A@#S2dWZQdOZeAY@c-;0+VOC1^V4T<9CaS_+AQR^GK?H2Gb@(]
#1IF4e>f;LL.6[YOK@f+IaVD5Z[g@@CPW8X@_4Dfa^IcZ;6CPT8RH:_F+<R9&9e@
PU[cOH=9-b^32V?eKQ]YVX+/B<RV,)&CVAE4G9e7VeB)8OM0e5S-DWXJ:V=bK@[(
\,I(Z9V0.6[a&RB#9PTZ+,gG^B0=1ZKNL:M<C6a?+-TI#RaA[_FA[d-d2B5eaSO1
,#_=4=+\32SN8BXbT6cSPC@2)F8M.(9_LcCa]Y=aA/f&PN(P6-YRJAL?/DCJ+<<A
38UWZ;VW#->Z[^UG6a\;0b#LE3=dA#CObB@F[C5FU[XEcf#9Vb/Ta7bUH1?CV=JD
ZP<<+3e;+FG(_W)MH1E1@5#L2$
`endprotected
