
// `include "../00_TESTBED/pseudo_DRAM.sv"
`include "Usertype.sv"

`define TOTAL_PATNUM  1000
`define SEEDS 100
`define cycle_time 15.0

program automatic PATTERN(input clk, INF.PATTERN inf);

`protected
\,>9/6Y-6GSg+M03Gc=TE&IM3RYP=10Ed:#]-EGe.TT0ESZI]_1Q2)bCK]^X-I_9
E&YZL<O/R#B^IR>#(R/T5PD\+c0Ea,8;PK[?,0):g<c-\gZa)>)8_-<:W717E\?c
:T;#J:@BTB9Eff7/@1(84)KSdB)f@FS^>_4CG]R49U7bdRKC:)Oa:bN&=4@H9d3@
d&9.0R<-?R_C]T901gBUVfMO)CSQL(9<\,IV_S+b;\VS3Z37\.G@\9(,8B?G\f6T
[9gYGf.NHY:UMH#;<HT15Xc[@#RGW7&I1WZIR#X@NIW>UZ(_4UYI;2g[\)?0X[K4
F1EM^<HJ;4cPb]gaNB:&ND@FK?JVCXGCG9E3aS<H51?e8T?/.58(50f8-S?6B@_^
VI1#:A/??ZfXf#W.2:c<W@a)SY02JU[IcGPV=Q]V,S[7,DY-2XZ6XN-[PE+_WOC3
fdPL0WN(HL&/[/F]@?L194O3M]fH66(^SX&68OZf>(LJ7Yd(aB@+Hg#FYUf,X2Y.
4dS0Kffd-JYF(+79F.eSAa\W4d+_TSZ<Lb#YR?aIcS7J5]\H@N81H<:#E,@b?>IF
CHVN)C2N]LR?&5dDP<+9b[K#I^4GO_YFZ2Ha\TC1@d0bO6XV]-,QB<@SgTSB63FX
QS02E9LFMKCLQ8U0=@F5[5:2-9=0Uf2bgIJANS&\RA?,Ve]9&YY^<;f=L^(<HXZ6
7M:aRP-R)-&<OED^B>\?0425Kf0RL.0V1+?X2NbLEcQA03;YTI=WPYWI)]LJDXGg
eTMR=86=?4E#eJ1VVFWXc9/[E@8RJ(&b&)W:DMDZ.6aR7A;V\VHP8Rd^1A[Ke411
4>0WYRJ5CdNEM.Fc.5I1J5@4f7aFL&0+d/HNEdV+d54Y1:<df2c/Pf&9Z=&NI,>;
c@W6Q@\Z/WG(c_1U12c:,+Y;NY-(cN1LbNHN],O>,aH7FA_<KE:&bGA(L\R?,a>-
1F,^WF/U#^)->JdMO2PKAK&4WagS]MDA9:TAA;<H-02\5JaYKKFbd+S0d:L^V8&T
;SF#Z(Z;(;9J69@\DC,Ie60-6a<5BG2fYNCSAG676MBQ8;@d6XUF4BH;d[JA#+O^
3B.[-Ka.I_N.@F,X8(\B?V1P=:A;M]^4?::Z=6=N61(.XEC[cU:=)fN:+J\(D-c6
ONXQ6)+J:Q&eG+g3W;>d&?\J0.U+dG+4G^3@c)(WG4WBY+7-/f#f&f.)LNDd5ZIV
5[T;1N7JT#I57UG;?H7?FYA>3+ZXRY2SR\X?FPM;;#0g/eT=-P1[S-:D@NMS/V,4
GSX;\?#)_YcAN7CA0AEPQ.W/I5eTDU<@:]?DY^bE,?(F/GZ5]/I(01KaV(QZ?fHM
f:f-[^HbF#C^-2X>5^?NY2G\)DX/-LEY/7C10J:<MBNaLQ:Q/.Pc1=HMa_,eLLDK
/3B#[A8\JT?#O7]<0J:dF4O2,AD9K939SJdI6VHX<JJQF9)QT/HMYF/CgGcP+4\(
N==X:^32GUJc_Og#-(ZEAYL.JbL>T1EZ+gXG2TFNEK73WabCRdL7>e6M-X8O<O8d
SX</N)LYEON(Be)M15M.6M(aPG9Aa])#NLB&IQG8R2fJQYO5(1LK6LPIBUJ5YcZc
QXX#R@bN&YORLT\K?XDB\<AF<PNBbd_E:V7S6R7.\&;&_bfc5MK2A?XZ?U6_[]O;
ZG@P=2??<<DFFF2fdd@)2G814>I.FaG2=7C/W3:c[)X?+PA^]3UEE?12g<UODAQa
M;1M.N^RHa9.,a<aWYR(,CGH+:?BS?>_7R)FL?+N<,--6-<JJdF5<[Z8YTK(5CXX
b<.4V3,RFKESd&A2;)O2X&=bBgP1AE.-048<(OO;:GJW09W:2E#LYG)_S9/B5U@I
>\J#Me0TF0PLa#<2BG9\G+U<VX>b;Z#YbHBWg2V\MVMAd]@/Y)HHV@YH=^A,:]PS
g#,@;,S]O8;/-#R05g#I+GWN=7^MK3e)baE?>^;YUL>0?I-QX#e840?52==IK5WS
@D17C@Z;=?IQP)2;N@F]RVY3&+gNU2/K^ZFJa87IU#fP@=<K>\b1F,WN(L.&;[4D
bL2>;,g;@ZVF/(XF;1&C4AHMg1R#K8E&70_;/3)B6\__6<X3ANQ/fG+SCKXe?I=/
>:4N-Wc4fAXTeNF@@GC7S2P1ed@&fZ#N.Qb76)d/Q>Z-R,F<,6^=/1T,21P35^._
A9_e[8BFc;_T6KcD?@/1a?N\gcF#-;@9TNT4^DTbL9<MOJ?;L867\beB8;].;c>d
3&c]B+8Z)+W5Z_Z@,KU36WGV@=de@P^6RIK@=WU6)R1:QPa_8]:)X8K_P7a;FWKU
FGGYIAA_-6SPHSWLb9dba?W^JDg-Y?R;Qg7@93QaRBOIQ@ULHH3>.-N&_+<1L5@_
Ra8f:]\a^[F@,]XD2#eW?/^7g6L2K)&NLO9#[FP70aG-PVVWT8IadK@D^VC?.e>^
E#W/<?RDK&Y^Z[Q&39]64K\fdO9,MWddb=,2:\^Ea+>7YEAS0Y/FF=915[e<cZ2+
a+8)L]g@[<)_12^\5LDgHM>LXP([/GFV8+^E@5e>\+1R-g8B0(EJ:Y0ed(U=GN[#
Q#PZU[@NOO<UHF]Z8VLS),d;]#8c:;b[gB9J:PQ^F0=VeIRN<Mb,e5_)H59IaIL8
(g9Y&5)a^QJ6+(YT6FPJ3GK=#6#W<Id__RW0Pf1W]Y<9#=L1NCbC_eFcX&]Paea?
J6e04bGS9EFX/Q\GF65[H9A&6D-g^GO-R/<e863,.4R=UC31]B9V\OTS<bM4-:,N
;QYB@:^g339(8;cOY]IHC,GH-(cGA<)/:M9M_LKDfT\X6Bb4IJYROXJJ&e.0DJB=
-#WFbQ#,UO9e,?Te1\f#N)O=^6a_a.:68e(7W3gMUI<eBR-MU&gMEM#S6-9Rf0>[
b9J>2b2/X2RW-cXQYL;.APfR#0.T:YMYI+SM(X;aM?K+B;A19B9[FK.HdFY,WYH[
],77OfIEM,UfKBWf7Nc7KV;[GY9aK]\8:BLgb-ALdLKD96Z(\M).42\GRG<:GS=[
g6dDgY-(e#L:UMR35_Y@&4YQZ=.dD>EKRL5gA#0>7.:\U=QPS<B9QTe4SGS;Pee=
^.(C_#Ce..(;/d0)402]]36JbM4eJ15UWO1.3+7W)0aFFD4Z#II^Rf<Z:2S@O/Q.
&DNO#.TXcT?fS+D/T)<(efdR/Q@fEe9M97JX_[P^cB&#^MCagC;+0eT(CE;FSG7H
R@&.BNQRR8?aa;R4[U-P=AC]_8I1EDW:#J+K:MY^DQc;L></B]BT.S)+b>SZJgTV
e#=8dP&98IFT&6:X1HZ&<_(0Ia8fB:LPMQ2.74CXU3W]cHgM1O3bYEI4F#8:;_P^
^34SRN:&d+OAgd2\GZA_\QBRAL)[,2TDO=[0^[&.0dM=-THH^TJ<&).F6ZN@Hc1K
EL;Uf&WKDOP<O5<#[8(:c;>0Z2IcXOFW+AgfR7W)5IO;/aTPP=7LP)5Y)DfQ@(Tg
:_K3,9-99TD34P1Z[4Q/dc6A3,T?M\+>fI+g.>fB2Gf/D7cI>V1:gPXg,V<J<^XZ
=8XG)5Y+2Y-9bd1.Y@1SbS.EY-2:Y2#HLb[b\I;Cf.B/@XM5B;)&VgD;YIb.g/E[
4Bb:[QGTZ\-g\C/LBQg/7+Q@89OA5?Y:dc?-_>A8W_X#IG;2DTdVOVf,O?Z1GV<?
HMI#2(eUf5ML;?]Kb/3HdJW3=DD@NC/XA[C>=b:5PS<C[Y=K)62BV@4UA:c^W/Md
C=57+^I1EWOCH7#)9SM//VSZgVEMCX(Md_?FBgI1U44PU2^OC(cB>X+#Qf+<,dbN
UEGI-,O#BS<UA@f:]9L8D9]HRKD(f6Sbc=U>P@2NZDXZU+U.)d-&>@Ae,fR>1J0G
a-94ZV\]:QY\^2#H1=,NM+Z)D&ZZO9_91/;?VD)d@\Za[P-@U4Q4Y<3RJ+aLJS(X
gLB,1f9bX0N<H<XW/+#a9;?Gc7&-G4^JYN[ef/_Z=e#47^F/4,GN&gf]59_[QJB-
>Y0ANDFWAZKSB#]NHO1Lg(L)/_4b3?_+4f\E+bZN+N#gC7Kb\,V+#SQQI/Y250>V
Sc4.8G,P-B:Q]F^Y-,&V;LUgZ=0;I7(+(1M[P2N,\SY1cIX47,\;BTdE^=1V89UH
]-#DdKdAZ3Tb0CC##ZgJ(b7LY<AW;Z0A-2A/2#OO=aQ&PU6WD/6\6eW;>V&ZJ(B+
MB5cAbb;8g9P1CAN?VfE5[PXEafM][3?YeUS7ec@F,7Od4G-9.G\+-+1E350Bg2W
_c_A<.?<++(/a3D11\K4QWR\MB^823702c_(,N2,/;<H5.SW)4U=XAca3:3&P^dB
,<<+LQeG(Z)HIBOO(V[MGOR.a0IFTe)-8Y;9U3@5bAV<e)ATNHD69JUD8I=A25L\
bB&4RWDgNca@f0D9,g3Gf)L)7@GJ7QKgB[W#+D:T--Z4G/Z60;c;AIeG@>^PD9(3
4J.5>Lbe#:Hd#N>KJePDXe6@Y.b\J+S75&3T?.I[\1VaOFE-Y@f/2CAU9<ZLGJ_R
]gZA+9gd).F@EMLA14S4J)@cYa.bYPJbQW#HHW&3K;?E2]>);W>Gc=G&E<FE9?TW
2RS<ac6MV-G:WcC2L[A0/.?WX1g3T8SI-f/22O8@T4/g3BCJO>@83).K4M-J#<IF
g)+.;_<)cP)1gA1gb=eP=FdAXZ.W#R0A._Y(=<HCKK9>+e0=I<T8V&>PA7XA@9,Z
L&Y0MGgIY0I<3;#VSUa89LS>.?G]=H=d=RA)HTNb/A@/TU.0UUHW^F(]2RJA06M_
Z8:2E.]57<FC7T?DagQKLUWLPLKR2FLE[U&b,26.U+<MFD+[2K8T(-Ya,T5-2?4c
26^Cb/K/K5)?0fI>^.T_5DS#VR0Of06-/XW]Bf[<L@&FM?VU3=K[b?L942>5ZDF,
a0]\G=9aVZHb36[>Od+_8d#;\TcJLKcX=f,CcbBc3aP-1N#-.e8Z&J7b)\-Nd89^
6/H(-30[a6K#<C/>>Y^S/VG/6Qc0WYcf8L23]XFC]R<;EX=+G0<[.QP_W.F@W,YY
8aeHCT]#E</.85QYBMF@/.=>:5D]A([E9KO3G/+XL8S>=N:_c4&#>DEY=+a[SD7?
7H]ZgI3T6Ka_aZBT_EHJcRM,&Gf+<g3<1Tcb7L.32#Vf10;0D<5T@5I/[<PH]]Y5
F[F3@:BIW0V3e=&JR)\g,bcF<-Y1ZO0@0U#FDSSA<0@IAJCASA3I#-5>?XL-WH&6
#0H7ZdWH/7QC7.T#G\7K3O6=\Ac;dMa643@F)2g2c,&(1Ke/LYJ<^HF^8TB;L(XY
O;O8b^12c\1XHL44\#&JI3J@O/NEXaOLGN8S\,)IP?bG-EW]J(ISg2AF\Z8J6gKX
.O_GDFSKD9P::2<BJ0#UD39+T4D-7gCY3H2-N(=fe)cJG,EG,b>&TV3O9gCNW?GV
\gRI@b/VJ#HAdW5b1U?@Z.WQa26[M-8&S]4.#UJT3/>:(2I&WO#.IC[/=M\d-XJJ
7L[Xc4;^UV:8=RUg8#?V)RD>_fb4b];7I4;?eFC@]9gg(#Q+0Z#5V3>CG2_7=6b#
CN#7Ge<^7L5cA8dHQ,NRP[T5dDVW:bLKb^GJA6=MR87b#&:FX0G/J+2QV9,51WGN
YEVf+\HPKDcWe9-@C@E]O[>F.MT9KU#0aSfI-M;LL@3EdF7-eDD9T8&Z83HcS-2G
?XHW#8JID=N3H1G/P8Dg4M43YQ\YD/2YP(7D)aV:g:Eg4ZGC<))[KHE]c2@K(ZYI
O&3<&(a5bYTTf=)Y#ab:6N=YEFaY?\6/)dfEc/eE522SL-Q-0P\\M8P+Y^3JP_I3
?,F]VQUe5?2QLPZ6<1O73LNV8:E]PXU>&65YI;#]UTGNgF^=QU^We&Q^b#]V<<d#
CWTPM(IC1>M,.]e^fO/#4HT/_E_BeBYbZ_8[7W5Kf>\.22e^8a3C>\HWd=S,+L])
.+G_UH2&ZeU@@WC/>3.-WC[=K<[PCEb,U@a&RQ3/1+,1aYYH&&a0^dN+CNcA9D0^
e35EeZ<Bg)5(,/?Ac1MdP??KFIJSD/LbY&:.LRY;9Y>14JXU:)_cYP7G.@GbI2,f
H]ed#479c60Z>K;0T7V4IK7e=egd/W&Z9E-6fRX_KU]S(Xe7C@bMH_:FKV\5dgAB
UAR-T1R]Y2I&DIOU0b5S,_<0(#9VRcD]&?C(2S_F5H?V.Y&,2);8H_)NdC<@-.Ff
;GZB<9<7AMGG>F@?g1-WQ5e]O.T_X731X>EN(C?HTRfg=gF3A2X9b,6C]Ha1WL/[
FT2\fPfW1FQ8>C3,d>#C47d26VFPTPgQ.aZEUf-GgZPbC9IQJ_YDE;:ZP]Kf5?^3
B+]#Q3C_GX#c8(,U-KbX;^DR+#_L8AS7_LFa(Te]#gQK9J-+X#PVaC?Zgb)bHB1Q
7O&?>OU\a#A8OIRPHH=5CC#8d;=cXA)QA[:,U<F:HfMf?LGVf]_0WNef0X[#fe?a
P0BV+5aTB,0<NCJ;CS_=Kb9F@2?[^VcC9),af\a[&_B>b:M3HN:C;VUNe?gJL=B/
=IDCV-6+7Cd6dT:&P6AJ5,K??1T[Y8;8]\UM_gD:N67?g;\FGdF7OdC/b0.I(FUb
84dVSQ3B?[YU9>;.:,92Zf?5c#&72R\fP+0\K=^EI[a=g&^1]M(@;UURMHKK.W)6
HHQ:B7ZeOTfQ4-NL_H.+P#)E)[N:V8Z:9DQFbCU)?YAOf=I^0RM>ZSHcSYS?_-52
KW3&Z[^O-_3E<+[=52<=a9)02;3\V5]&5^QRID_ScEQ)NK?]QGb28J^?X/f&eKZU
K#P93gae=TN0dN[MRP(9H,G?9??+X_#F(>>\)QA<&X8c,CMDP08:7?9&T#SbY)-<
X1E31UR.c4(>I.f<9?A5V/WS(6403O>KUZ@-A8I/P;RRMUYYR1ZTPDe11=bI_@[Z
-ZKJMOd6U8T&>W9LTcB5/>GP]@J=?I0@)&(NSIEBE8=K5O&6IK.;:4:,P1=B5#B7
d.5LY&JP8,GR9=CK-E/2Z)c9W&gE5L?GXXK8\G&3T9==<f?S_U0=E05#+H_fb<Q8
_3;LQCN#.92Tf;FO7/Oa-eV-\KeCXO<ND+>AL_68OfVb<7-&65\cG5FNg/]279=Q
T=+Sf9O>Xe/d=b8/NH..M??RIg8HPO_J6gJW];U&Vb7f8\WN\7c0K>=^L0cGb?PW
1CFS9E\ga/MW1AN19IUT,NM>dgd&AeT-OL+IMf7V0.:KI/EMXg(AW=(3:9X^K-b?
GCfg:NfL\9TTc;>_d_.G7b7(AZb4cb(6f3MQ+1[RdYI-,UHM+W9HW3N56L=YH_J?
5[bBVMC>GF.G1F[EF@.?.3/QV6cT/PUIX4V+DA05DBOG.bN+BJY^<=SM6JHX9X@=
6<:cJ1K-,e45eD3L2877.[Q&DWada:C.Q2-=P2a;^=(F#\ED]6H_1[<\<HQe)/P1
9P+PD5-GI)d-.LAY.WGY\_(X;:I3#a(Y+YON.ab,JPa@NI_K3U,@5K7Pd\KA(4>a
K2G;L&+D.KSPUMI0VQKX9+;0[[).N)-R_KM.5HEMHD5dKD2(?G0]\3EGa5_L_39L
:__,E<^541VNVLdH6W0\>_0f7+;e+-,&CV@A0AFLLaB)0g+8GKbHZX>0^XHb16bW
9DdR@>dOZ8J1d<Z6ZJ[gL=3+:62>FE^HJV-?9[:4OR.4+AM<Z?#L-J-LJ33dd^&J
P>?5JMeO4E-FUS+VUXa[6VHGHL37^_S^PT-eB@18RN<G86\<a(.=:,2P][1(YHJ<
>Q&eB<JWfWT9N79c(DHU@2c=#8IWSG]._IM\fJ>&H1F]J6E&]1+^/OfgVOE791X#
gc@#[a>NAI9A&39g=F+XK0c9MOI8/Z_O-XW9\>YN#Z(;D#UaJ-OJ#K<>fSGS26_Z
U;2UVef=519&8JE(#0[.<\AF-)8CRS(=Uc[+<PP[Q\H@(HfLG<W5HKG(L(QN++2/
V-D:BDX5647I>IWFdB>F[RUX#&UDEeU^=2E8Z_e[Mc[e#?c3ef2;RHQba@Q_@+^&
M@]1C(NU0D20NULF/9f1#0__BcZV@P7#c6.&N0I5EIER:.#dC2EI@8PKE?@@VLOS
WYN#^44P.K4F/)?=NW#5,aa8+,2]UCUP-g-dgVcD>O/O;_a;[M.+1H64)]f;[)&I
22,XW]EfOX[J\P/J\Q&WM2TZ]V6BVUMg/c^2PI-IFTJ&SeUMYY#YXOJ4;A[3VYM1
EI8#\<U;=&ZCV6^\IKTfV+^N5W#D1Ae5ZTSb]HT64K.38:@+->A+)HT\P1Le?EA_
B\S&>Ee1SQ4YW:_5Z>e7[L6654Y5QCR.]fCJWd,2X(e283.ZMDN+6cNG0TW>UW<:
#^.FHIZJ@XML4;(4ZXV=BVP-H0=gZ0P7Q;c\S>=M(f/S[C\c5B\N>Ya:#]6EE0S=
>P>JJPFX()^XHDEFR/@RU)=\(5G0=_TFRaHU^Kd^KU#-T,6;/E[9cSACdRH2(B5?
=Y:TD\C[AOX/g0Q=Y,1b](-=Ya?Ifdf6:0+^LS1W8CY7]M)7LW76@)#[P1\b-;g.
)@dZaUN9?W\:D-T;.M2bF/aF&YK@>e4;T(]30UgPB0\:<Z[@7G<+8<4Md.:L>-;Y
]g&NUSIMRAW.V_Mf/W\Md65Q)0MC.KKP7c\(?fFX<5IDg2769[1ZaAYfYXbGKN(.
4DA/77LWdV6]\2XA+AD6+g>-(XaJ3__PG@.[9NFSb?_NF8fX>L,12.>Y5R<gIAG)
/f2C\_2BAY3E5#aVTA-3Ad,W)5)@=:&4gXOR35:KgG9EQ,K;/g2QA3M/gIMI^;cf
:\2Q0MIX<,B8_]WY>7Y-g1.b.@35(Z/=JO18PH7<@BIUB7=3gVdeA^,RX<4>\>1/
V:Qb74XCd-P7fF]c+W+T-BK5/f/OBP&^E)D52b\KLT)Td_ELCXXca&,3C,P\JXD&
N9RGLY]MV05?g,+7&O#ebC4cJJMfH=J7eGBJb;PEIWMPCaR9DBM-HaH=G3<2SE[0
A8FJc\V)I\A0P#(EJPT/T+d].QU-geI^>O+b2bF(?OSY<_Ua444AQL@T=:/5\Z4_
&C-a<)G@N5]&EZ7\eRSXcTF)WG5)(O-Xd/K:H61NCUH.Id/.?\/;<-7QdGF&7DDT
D?)Xd#2@<39)+JZM4RaYS6I2\[#RbEM^&PE61PVPEe.fO1]]9c.C>Q_ZD\OG;2S7
g33RRDQ(+[7BVZdKHXR^00K74b7e_aO_SgXMF=,5:.f4><d\CXOXb<9UFJF2;f]N
ZQU&7MTVCJ2F,f7NdL3VDGC0-/ZIAb:US\Q&&e-&(@AZ5=eIQ8LXB)#QVA1O,VN#
3O^OJeK0W0OQM7Acd;deFM&&E4]POALZITW7ICODd\Lg.EDGTLSYaHS,NL/&BE^d
CL(=XLb,O]JDGdMV[JBA-_dV&(0Pcd_<[R(N-Tc^X_]MO1YI\]4a2BJ+a([7D39U
)&,Xg_C]YaSZdRIG60/F:(B#Y[6XY[GALf4GD_,BJ-f>G,0A>#9aM]QN-F5YKJSa
Oa8P&XB\QVGI<VeB)K^R8@d]_/AM]2/<Z(E.>R]dJX]157I3=+>2]5VD+9<6@0f,
>,2@-#S<^A;bXKc(F,e?60IdQ#O:\&MWLV39TU61C16(ffEO3bKY<;(AN8OS9U\>
b]cVbT(5[P1\2^LB7GN@O82.8+3HE^UYXRgaA_?]XAB0;TgZ6Oa-N\)M@fRX>df+
I)9E-D<[^)eG5IUJ&?#WeZKE)V]R??N8MQANO:KNI5(NJ?a]W2@?5#+W:V_e4YOd
(H@a^K^fAb\YSa6We(&#0=cAgE4Qg1d?2S-SL[5427:PKI:^87-8##NH2BE<BA8.
_&XS=BZ(L32KcKEgc7Oe,b1d4ZT@H.,:92WA<(+10,gg?@cS4MC3c^>_::4fVN/G
UI#.<15]<P6?fO34)5VcU_44_0#0fRJSOb+dJM:R[AHK^G231^WTP(aQDb\ILB37
b/W9eQHTgWX=f^-E81B,9Y&-.K@=Q8U1LZA?I,679BcdR..L=Y=2P882LKD^eQ(\
[a;^eGeRX<;ZBO(S?fKbHbU5dK8/RRW)adRfBK0R\Ud+K#I)AZ-PAa)T#_LfTfd;
TOeYM:73J0?\E0I56=>_]?,76UD7M)/0De+1,P)(V^d)B?=g;@[]a9W4G;(N41;d
O+#H_dGHEb-H:dE]R[:B(^(2)0<&NYMIa9.I_7YWR7+<bD;VP#;I28NP66#H[FNZ
aZ2EJG+f&=Z;[#=#a7OC.CC-f@GTL&c&D:&?Q,0OYg]<>#E#7K^:SJb_/f-JXN@X
60:M1YTG9Z(a6aKWLTa3D,-dNNY?,5,FE@M<(,C:4,Oe>[FbCLY[4==A:dOAAWd-
:Xg<d0(G?cRWP,NG/[NE=3L?b7Y&LL6SN+^#5^?FTDZ]PbP:IY4@#<f.c]9fH469
Jc@\b?3[OKU13S-,Afg=ACIP2H0IHR?4g7RfQ6&6^,5(Q\[XMR^)(76@4;-[#Q;d
S1;T/&.5fDd3]<b:/0(:,4TUR,[YCN#IeG>Nc,LJ19_<T0S]K)WQQ8V0./GA?C.&
W0;g)c?f]aOMa)31EgR>>9=#VeM])I]/S/EGK62TRLE3[M99\b&De)G5&#>4;OBI
VYYR1@X1P81D\8N:+ZeZ2?&#g6X1\#[B8KcRZ>gVMQWQ9WK8aY2.6B?P7JacW6S3
(2^F187D\fdQT#cHAG_X;)<.T9YW+fOP^?gf7T8(6a(/7NAJD_6JR,aCH0@Wa5g:
\G5F;gSKed6VDF^P,L@)<>?3:K+0(_W>[BS(2OELd#\.6F;8?:;[OJbCN8UZ3)V/
b]D8=3GK)=faFGf,+EG[9@JWU2\N(1ZWFQ8^[=IP<^D<V.F;X-M&)^X:PZL]G\UQ
[eRBR5>#CS](ORN(+C6:^A79Wa-:/P;K2ZF<J.S>QQEDO?IT#XR=LJ:,N@K=M;<Q
Z4K>^TFg/-[Ma&&8Z?6&S20fI5dX#.d\GNC:JFH/4dPJA+1g-92)C0X89,,9fNS8
39ANUF+C=RUAOX1M]PQ0FS36&3YQA5Ha,gdP#44D6VP/)NQRc4b3Z107QCU)?Ya&
E=RR,cS64(C&_S2YWf_Y]92JdA.;1]>Q3:&9f)cIN?A8-(MA#gM5.T]6M)LOO5^L
^e@EM#8f?8bT)5gS8)572]G3G\JX;&BR#DcL7X_I=B<B<UW1RPaM@RXe&N9NA^DE
(XaGRgEA50Y0]_&[fOCHP&?-K+?a@).N1M#QG&E4D_[5cUQaXLHUJL0a6D.>Q.34
+D;e&fbTdc=>@?+EMDDUET3F6FfVFY,UKZKfQLD4QfILa:L?UH-dR<_g=G]2&fg3
<CXA^Pcf+T6,L-Q:<4LNQ<XU:P3C8/AEZgTA/0F>P9@b.b)V5/6P]+AE(YJL]PA0
0E-M>BY75^-PS1dfPYbLb0Y,\f36A?/cRb:]a7MbYY20\TYc:Y<4,fGUNLc[8/@6
UPa(CX#QA>H&)5?Y,LK3HJSI3A]-&-OS?5G1L4CTW9SBQaJ=Oc]JBARGC>cJ1_AJ
#/bRHgP(Q2.M]@3V+?8+5)&]/_H\>/JMa]:N2+NJ@dLZ,G1..:P1F0O8E\U-XfKD
M1B8fJXF1(e:LT1b?IgM3cWbQCO6UdNZ3DfT_000T)HZ4,Y[W^;+_T5D.><Z&^FO
2aH#+;b@^9M5A:B&8I.G/&cERg13AF;A@a6c/2M4PWWH+.f;8gC,-0)bc\I2,-c@
P(QSfVgabTP5YLB)?&)2<VLZ+PC?:(UY),eQZS+/;TFT_,/J<If^,R:0XG[+LTP8
PA>LJF=;NCggb;+daE6J^Y9MLQ\8N^_3fAag867g)JE/9SfQfTPSD+g)cH&_M_c?
BQ6>@/>EV=S[?O#<SE^5&),^\7PS_4T<2@JaO&a>&UI47&8Q<a::M5dO##R^GJ9K
)7B@-QJf:;=K?VOf3Z=FKbcT3bTC8A&6MCCTP]YZ>6:Ee,>/).K,.)FVX.HeP>MK
a56DTUaOMJ66@gcLY1,&#GIH2Y2EH>.GT8DXZ#A^>^f4OFW-D?521]F=+I.I<MF?
MA.[LS)XcVW2?QUQ.M^Y0cQ3^)G@:4Z.DBZ.bGfXP/ND&TK0bYYc8KL7^-7<M(N5
EN+W&=A<CJPV,;C#P5#[ebcF/dZPDEb??@f=[[.>2feI3d-N_V77dO+=3.)]?.60
YDD_RLJcSEIWS6()NZ&:OAD<Q(P2TEFSc9VX6c6F801\C)J[^9^)ag>#_4VNM1.K
G\bB;H638_D2gAAeG_JI[-TP1G>(D0bgTG;,R)7&W^U[I4JINKI(]3V)FEMYK[fg
T9(KV-M^@549E->DCO>&V75QYVIH+S_-=G.50C23,dB9-5J>69&/+E\05\N]9^XI
Of)-Q0Xf3IbaQHO-IE8V=b<Q,N@?dCD;:_PWMIfK>^IY..aJcHeD=H[FL?.0<CEF
TE>g],0/7Be@;+\\>1GUB>60.U;U>8)),]._X3fY5C@2=Gc7_(^]552V/9UMJRE.
.M\NJIW6UB5_4&@Ee0R\Dc(8G:e&b::->&d5B4&JgWZB:;1P74W+Ue)>NXK2@LgF
IdTa0U,7P^e.)^S<P:<@<N2)BP[YW]I^@<I1/TU//V4/ZM[g/MDcBI<CW0+TLB5#
(=&6I74/>e:&\3XXaId@f_=701AS\N@8P6;6>E7;M(I@>gJS3aSccQA(GTH_d=93
\@DYK^W]&a]\IPGOb0)07AaO@aDH@YKYVK4ACBaWC)..?2(WN:DW+K@:3Z>.5dB+
5KN8ND10c;0G@M,;#G8[JESeDEffOPLZNMNRef-(ML:3Z<,L;:,9H+&(?f:AC:D.
gT8=;EH89:b=#>e9ZZf78c76(d424W6A2B4LSe]>=HNb0P,(+:8B<<2&G@Z<FO\<
-D2,5L]-?AI]D0AdfK[G)?.IYDN/F4[EgSR]bX9D>,?Ve;6(I>J6X4D:>7d9+2K?
[3CSWEJ]TS6XC7UX92@?T]UZ3f2?E8-XT46JZbZ6:\MNSP=4@^5FX2ad<+)VQH0c
R/UE2]H2)JUe&E=f3TJ1LPQ]Q4a16GYg-8PDS^,:MLRZM/4?OE2:(HaZDL[,dWX+
3gT]OdCV]A+=d;A@?+D;++c8]T?L=^A_O4/9?SXc_=NCH]H)P1&&]:bbKO0eI<EC
5Z#S\0)/aDQPDcS353NM71#:LBCKD/7e[YE5fd,U=:Z5(O)V6&g<@>UHd<=?R6-f
W\&SQ;1:)C>XN:9a4O(N;GB3[?C3Ff1K@3RfA48PX)&,JHT?d>1@4)Z:Kbc2&)LO
8A[;]FDW1QR\\V05GQOaM9gg]Y;1ID?TJX:IPIN0c.X(/g->b3I9?G@D(CFC561b
F+8Ha&R5E+/IM;c1gF;?P4:Le?,>+cX3WDe(U+I\BeD=YUB)>E-Rc5@75:(f@)KD
IFU:c_KI._3^<&=aJ.NVEJ^5L>14().@64MAQ0\[,0^.PLC\.B95eF6aDSb-?)Od
/6H&EDM)?;;e&IO;;;YZI1Y(eOU4&K4+-_5TRG4e_FXIZ8C2dcd9V^+,HYRQE\._
J-QJg,^e;RXg#=;2S-X0g0NX3_&UNG&&O&<^9?feSS11X<9?[.2TaP;/SW/B4/24
Mb9Kg+A_X6FNMOLBFd/d8)=;\0)17&JdR:M2+8?Ze2XLQV-f<D_44MJ,B8TVX(V1
GX<Q.g9_:BXg55C)-?XP:U;e2Z<cHIbQ)Z8A^^UX<HA,E_(ESfYd-40R/^CGY1]]
KZV8\&IJM1@9[(>VF_^OUV8/ZT9=gPQG\4g8d9V4&83O+NBdGQT3:DMaF4XV82/U
P9VIDD5C\+^[-I5X>]R(&If<9Z]2F)e\1-(G;c&]_+fJ:>[fC5fS.\;ATfcY4ID8
5\87QQ:V,4_:2QKg]::<B-&Z^B4M8W#U+1];OO&QN+92IH?&=M)#b&CX^+ZOH\59
?g[X;A;KJ;eV=4Xf2MU[?e9-0JdYJ]BV2QTc3Vg7UGM)3Ie0EM+?+FJU2Z._KHND
e/g<gVDg(H8.d#6ad@OI^]R+bCR:MQb)I#FHMTM?MLFSQaA@LQ=>f=,KQWG_Q8QC
<Z_CNdVR/JZ(aO\JaP4EGX7eFK-,d7DM8_YObe35]3a-.JXg2Pc-]F^L/PVKg,\Z
ZXc/8bG,_AEX@ZDe0fX=[XF6(K4&NR-PJ?H=,8_gWF/(bA?TM/QUCM.ASd2TZ(cY
C0)PO.63g.C;L]fZJN_?O)H5:>gcCe<T,+5T_@Y0[.V9YJ@ddL6DFPF:7f=,Z>6&
+dR1=2<c+dYd>^C8f5:0IRKY=M@0=I6X#C.WaD7=>.),cFfIIJX.D_]JG5I+JeTN
U:D(IO:OYb03LD6XENHKA?31&PE_VG_3YW=;K2?T3XXCdT399PZHMNY<_gH[2JO;
3P>V]8O?fRc#g.7-1?.RgMNANLA]T;Z9F+g:+:#YVL[I+MK,J#M_QeU)NS1N<&H8
-@G6>QS2ZaW>S8bIaXb+5O7394X+[YE+)WY>GCDd2We(?_baBGSgATNLILG@SGLN
X1H&<Z9[U-,gH:Cc&^7Z:2(Y,KU4\ea<VQd\C.Y2CIb51Oa\Eg&Ra_J//G/\(BTc
)G2Tg#Z<M^;7E5QQ_=GWSfJ=d\0fCS0BB>_gJH8^,>W9>:OE?SS;;[EVffA;WIZE
P=HAQA/Gg76TfQa6POg2BCd0J?Se0<KWV#LRIWX4;&1Ia@S;&_3N95,SCU(FH8LL
RdE>_3Oa5OWa3OS7081T+8X[_c]ga2TY5XG>7FgEPLYWH(DT_WGDXN.)f@c3V+WB
@.aTe8KSIW4H,U]AL&TgT<74JEH.&Ga@5B7@I[]JPM/0@B;1/A/JF+/8)E3X[;2[
.UUXT15W^XGYe(#NJH:4+3_7:\0[>RPa&4:,P-a/Pbc.?8?&7T<?)_QT1[VXa)Yg
JKC?Z]eV3^0;9VJ\Z=VS.I94\XA5<SJf0_M/A\#M.&\;#Ic;6V]5aG9,T=\P2+-T
3fJ(;.84[?&LCY:N),SCbOM955K<CPFHfgg55_KW@?<[;g,=8)7&6af9HM_^92UI
84(&CX<GeY0Q&2Gg\KTf[N5FbG7Y)#&/ca-(b2U(/,?I7[e)a=g7,-C8R3M2g0Fe
NFBRI2W@Q8J]L]e=4Y3&4?V1PHZa\EU)LG9JYAYMgW;-fH(+(JV_8XX+\TcJB-Q]
&EC0Qf4MKJFBJa&6?YCAZa/S)(4bG_[@6;Q-ZHWg=Sc@#]>LbZN0_f^?FfSa5f<2
dc08GQ2f047<V&?@1D>N42C<a/(HH0(d608Na_4[F^bEK/6d;--M7V/<SgOO]Ub0
U19;F0T)N#NWC_4e#1;.(TDT=(<dY;b>(5+#KV_1E5]W=>:YI_>)(Qa5MIR\9=X9
YR:EfVaI[-8UGFD[971(/9:D0GC63_OMN:Q4fc06<8XQS[J#,.c1a++SXHT&+Y=H
AJN6DgH+&Q;ef0N(dGQCTCPcRD.#bT<<BBL;<A)-)1J6.U<]dBQ-0@Y38W.N2+G,
8f0[dSN^4>PMAY7,M.bgD<&2,d_/a#IDHU@WZ:^,3<T=;aU5+48KH/G=M94cQ^6Z
;+2F[R,._T,YN3P(QQ#K1.<;&;L@b3WL;SSf9K4#XR2Ba(T:C+[:5TVVZI7WXe^.
^>SS+]f4+/aXXef)&3+^Q5[4UI66L>_A0EZ5IO#^#468DFCc5U)6BbBc:A@8>@fR
6:Q7(W,UCHF>F#P5?TWGcE(?\/d+9W.9I(L5aH];^VLEO6I42Lba(\\2Q,NFU[c>
RJ#E;ZVA.PabR65TL#_LOAOKKO@2b+@LFCaZ>b7:[<cU7bUT16HaP[E4S)gIYZNZ
=F+_[.SBW[b9XBN)/PF/B3&_/+W7G6eF9IS?#Y2MDf;-BO99BP1^4N\XZGE,#e/P
VU7XN-:?F+GCJ[3[-U(/-L8X;bIaP6X_f>_XbPU,>W1:_W2[)c?/RS^=;KR5I?&A
Yf_9HSH->_<YYZfb(a3K_b\&R3SBR?/Ye61OIEMa[F9]1:gX3BJB88NLRU:0LA7Q
)FI53=eJVC,5-<dB.YES2E@U.ReQ5-&eQ.@0WX_@Qc/7MAG]3^VZ/1.<)FU5Hd=)
I=#AdNWH\eB(Ab9V9&@(U+e^,EZ--Y.S=)M4>\/Tf?H;.DW_DSVDJ9CAQZKE\LU1
C2^@<fdB<Ga@[^J78&#0=Z[Y247X\1R0AH,OYZ<X-,AB1F@P0(7RTU#PWD)QBF&U
^a(+J#1,15e7Mg/K\U=9V3M8<f@M6.eKZfBE+J/P185FX4YT<E_M6.FY1fGcFJ]S
(]:eI(:CQg>SXO[@.;7G=d]UR&I/L^RM5X5-;7ASQ\_eV(@]>.Ug-SCcWR)LP:G=
7L:22NYX3_M,TDU^/6[NBTP4G?H5&XgS:1UKc0(AU2XaT4^_e.HCMW8&[V+3OLF/
6+STON-X.V1C@U6^c/D-HI(7ea<?D5_?eJW?^RD:Cc[SOD[O7NIH,ISGTDJ\B&[E
1YYO1).Ce(P_7ba[TTg#^E2W&5/A?-1^HVDX5aaC&[1L>cM?6),6-&AANaHNDTFJ
^SM5SbadVUe.#JH]Y<Q?&f4bG,gd,I7d6WA2b_1N(R)@MYXd[_^EN)aVQ7<V4W+L
=[d>@AXWQDKQKQ\KPZ^1=f3S669#?6Gd(1R[[M8T[0dfS>MIY>)@1OMg#,FDXW.V
eTcIQcI4?\@aWWM,+dWPAT._HD09;]c^_-:]#I^>WA]^DdS_>gZ74/SV2F^=,>+O
-TT#P9[>_13/#L/?d-U(gH0BRX6LS_FEEeJ)AJ2RG27CLFJg<_)U6UU\KJNOZX.7
CdZV#-J(8A/gL)1J?AaYFR4VcD@0[HDHQ0DXGMEO-F:0S8I;6TU=A=DdS9XH5,HL
M(QJe>#aBI>cM9+DQ[-3e[<O9P1;Ye+_OUE,6I?HT@FG_5DC(1OS7NCaE<58939P
,FXg0F(07Z3M+LULVUX&BfTeE#A:/RcBa+5RX#gPU\]/Y](8V&CA7[IT?EK+6P]e
FYGb/\^bLd(]0DRS,IDK4#3b(;W9JPOYTZg;PK@?,Q>NGU^-agOX^7M&GP@U@4+L
9G/ZCB&V)-(OgRF38V:)Tg@W0#V][b2Q.BNR.MVK8ebIJQ,(d^#]P//bN?SbI00L
;2JV0;J/FbM?:a(YT?V_@8CP)JgN]7ffX28<9c,GE,Q3Uc,/36]]9\@:-+9gT>d5
1\CJOK4O7X<[/HC.O3L^B2(EDbdHEFDOefF;/aR4XR3gXB]#=7A:.V59LPM6&0O,
R?EF^QaQ]dQF.(a[00P\2<#OfMYVIJb#TfQX27ELb(/RFad7b\@)DXgCP=RU9G?>
+/Y85PYVP+LLVb35>E-PN4[N0QD_2dS4bL(4Z[<ADC]C\4\IGFKa7]Y#9:<KJ2R4
VG69CY8P]aH>N4T,dCQ;7S:gcbe.Z1^Of:JL9Y&1XIC&T#cCPK?.HgU,/TN,(&=g
3e3?OS.ZSBV<O.G24U5.STM]4(H<>.^)gUX1FX11d=O7TF56ADR&^61fWB,@N&,#
MFIP=X/)-^FWV-^TA/WKP?Z=>_J3.bZQ;_G&.<eX2.\MD=1TQ4#+\BC]5a<RYc+X
G0JTH^Ld1<.UE>ZE2_-/=,/8E2>UJ4Z\&&g^I_OBK?YGH?a3/=aEfNN9;1V>&a3Q
H;SP))A>6YeIND83GQS#.0D[;K(,[K\66e\VcHJK?_;LOeQ3PX,L@C3cXN2e?AJ]
a708L],]V_1I<1gHTe94TU<KFU3(Fb89LU-I40QddJE&DM:(LdFdE#+7=KF[Qd([
,>Naa^WPdL2Z=KN(]0gX;M+<^SL4C#5INYL8Xa)/K:-\&H<7[>F4MX/UC][=EONR
)4d4NCcUG_KefF0EM4(G#&_e^OK<C/XYK1_-](D<:OXXQV=83,WD-eWG1L(,,fc_
7W)DPV5a8B.RbdcdF?Q&X^E?a86L4Q=65Y1/Q1f,NAXGFD<=<R(;EQTYgTbfN-^a
dB+Cg32>4e?aS(^I1QLEW,ENOd-N_T/QceH_JFS+P@eWe8)UZW4<=HT6GLC=Z\]_
-VJc-C91\/R/?N;J@ef-BD(O[Za/Ed?3[IWW@(g?D=7NR?YO1&QXE.==;,4+^AVM
8/A-2-GIOgWBbY/UDI+F^5b8eMc[1c=;)1J@JPba<cg_5aS/?EJE2c&44b?O#=3=
BBZ:0]Y0BR-\;[T58XWQQS_c]fU:Rec2RE=8RQSV6<:cU7Fge017+I]:+b4Y,eT]
[c.4_81-3CK&5bZF>O7(d<WNc=SOSfPO082<NL=SEP]:#)-d8W^]Lb2Y#ceba=][
ABAUH&=U[[:C+UA[_VfS)JCC#MB#QV7@._:/?aF#Fe;FL_F4\VX6LI8/1,:g_d(1
#C=/1Q-L1=dWJ1T/SFAH-X07eB).#LF#PGG)XgS[^;JTTa\9AYf0R6KgcVX[RF4J
#A,)\8.=]WQ2Xa\JZReC;C:RG>f36.LFMGUJ#/._HM80.,=ce&A947dF+/Qb7O_L
42\KO8:d-V0;SW(>W^0b/(>J)R>gV<Td@<Y9TG@=@3V3<ZBDJNO@BJOI+HLGE0UE
V5GYg,R:LeWfLR?_OA@BN9,=@a8K3+<^R)eM+Q8K@GQ<9_SO-Aa=9aW)4?[H,FJG
_aDK7EH34M;@H^H)26M5Q2)6Z<_F>7c.Y.AScKSe/-Qb#CJK9Xg7VD=4KU6b6P-&
KNUd:gW0ca74>+5JFeO5f^5;:c,(8bW[K=.BB4[X>ANRFOaHa9F\>X=6ILe\\aN4
1^7@7^X=8RgdUO[2)]S:d<_(9#FSHDA0H.gE.>5B,D;;V]#I=#AQWa(/Z@KBXO?f
T)(P1aAV6?F=<C1[@.Z1&^,)(#6R,X(aVe^g.@CI&@.5XA>2),2I1.EWG7Y>aB,&
E=X09RVK[8K.:\TEeF.SeN.@.&)b1PAD1Y1-GP;94?IOE3)ICG3GJU-Z?eZgB/(f
P(]HL27e]1M,:0@D>E5KW3edTUB7I(:K-JQ>AI^9^9LLZZ)Tc_JULKV192[^&8)L
\58YV\Xd@-?@U[1e:M.S&BYJ\36EC+3MKSWLX-A#HL(/L^Zb,16:d41;aM5FOSDT
CM(P)9/\)/J&?(VU8d2]e@R+.N&A]Z0b+T,N<7=Ke;;^Z;PK#827E(2_T/.;-L]Z
>5PEbHeY-G;1U4;K:HI:^^)Y9bZ,/_BK?BF,G:-LacP\KQ1>]HM.I831?gC@DN&;
X_<Q#YR;.(,](#?E4)8EFD[:c#8.Y#A\O@gEc\gR:H/QAOAC\101^2?b]=NFg89-
1@K3\=DaIO]1&E[/L&15:=D;CQ1T&ES#<K,+Z(.5^@[E\Neb3)EdC(:4+..DTDEO
W)>B)9:N(?.:MA6.b&7N[B-#D[_M?P1+8ac)/?C.-PRZ^(BebFaV5)#&PKUHSSC:
/20Dd@=,I&dI8D^I5^_L):MZ:SWBaCQ,+<Wg0C_\?FU]Y0Jd@M?2XKH6cH]S;V_L
UN6A^]Ag5Q:dd__]cQT<]K/+BVO)9ICC-f2Q[,4<C#>f9\;XL27.OVS=B@9EW^1,
@+K::cX1VKOAC[+fE?FNX>CTf1P\WY(<.>3ZM_(XNb#T8=Y;3,7P+ec7M;:d.0X;
Z,^S&Ne^DFDf41;OZCD39XE)SJ140K&aO^FBbLD0R78<_Cg3fQd]B3;6Z8;N\7b9
aDP)>?):eNR>O;KQ#Y@E)?dFZN).K0BdHNbfgQU58<d+C2QNKEEK5b0)GQOXA+6V
C?L5#JPWCLe=,#9bTfB(8GZYUV8Ya7A7K>be@/POYKYaLS)a=&WDP?d)FV@F(T.U
>0;HL144+MeJ2XBJ^M^73HTFA1bPe=Rd8V?#MLf.R_@(O-&/?44_,7Y.dTM@R[NP
^cB92a;e=M#G:WeD=>07\O:.[acW;8==FIcNMIYJMZOASRYQ>(IabP(XR&e545Q?
e.WW-NTDafZV:)\EKE;gFM,M=2OL2@e6,W^]<CM)S,>CKL?c@;=;?7UB];<KU5ZI
)]B[\WfWIG9X\]cX253e?I39>8M-_8e_+1HZd#1@Yag@T].N?4G?4aFY3RUB51RF
HV.Tg+2H>I0:UCR&9(DD+OZ0:/&+GL@JW@1LOaaU>/gK1HV6?/RP?]@SF:c<>H88
HC2W0L:A-O]URX/02JM]&G(G;bVMNAf;DN)8>AJcSWS5#VN[C&)UcgY>1)#XW5aH
0EX+T;UaHRc(dJ0&2(5J3))6;gOHE8H(9::,BD1&c9O0LcKW&A2MVH>\O,Le\W89
(NQ&#1(BgEHOFEQS:Q,WbZVAHefES?3U_T>8UA];T#ESAQ-F)H(U)ce;WHXfDN5g
LFT7;#VE14[]Z45JTfT58KE(,KTYZRNg>+SKQ?<[NbMf@U9b\J?TP5=3K:XHVHPS
D=g1LW&3)L>UWGFJ;LReO@^g:KZTF#V1\>Z21:T(G.:3DMD@,(4=F72^H2Z61ag^
1/HOOg.^J;f27^;IGZ]_J-Z=,\J+e.LPDVb;#P&EM6)#b]-\/>A^EGCWS\>>&IR&
@5A?PHa+ZXUEMZB0f@Je&b+R<V3B\dY8DW.eL4MPASWDT@-&CU+b,Ca(T3FgZGa[
A&O[E[@63PYaN9c2S;eBL^\QdQc#e@\4#K:BcZ:2Da2>M]WY+>eFJ]W\HM9gIFfL
FgbOCNJ1Sd;^^)POW&[^:2&.W9.:e00..dT?S?Y)Uf6W4<N+B<S,8G3_1J,,1e^9
V;[WP>JBGGXQa?e/]e-O1<S/#16YQIE7K]HQ:6_BRNfN.DC\P(B;P^FF,2cA8e<,
5d9#KI\/c-FN^=YfI6ZJb>AfB\\@e(;P7U<E)@gba=O9;-;[,3>c@&0^I/\9]O-I
fUP-0aGFO@\XEKcQWL9Q60aEJ3VEHI):X>eQ,?b@RPYf3eUZ=Q..]\[1ZRKWNLZN
RAM(Q41NS;?WbON3a-35I-f]AYCRf<B7TGIFgL;?KC6)3>RP3(OC?F0E7.X3fCG\
JY@39HaP]AF;GVe8aKC]@]6(JTb>bHJTeWPPU?/YcfAbH,J^OF+?C2?JD:QT_/EH
4Kg^U/^;g@)7+BB3^:A7@O?_UY::#(gfQV32:Y/4H.Pg7c>JS:-6O(^@5e&3=/8f
?Q0@)()E7#KFQSVG\VCOM.57.c;WINWV>Z>0F=N=25O4DgQ81_X9;^Z&159E4Y7L
]6[BM8\89b[F1K4TG#__)K:]+K:8C)PL(E?JMgJcQ<ZA_.)4<fc>f2F=EV\BdJOX
>H@+(M9_6W2G=T.;F9]@QBY>)g\G(C^)&IC?<\B547;SSaYWCV)f4]F^?9F4g47b
I<\2bS(R9Z(PC++K.5g\BTR=5EL3M[G&:<6>N-)Q@JOX9>5>0&f]OPN7e:.XTR4^
^gbCMWI\efNIa14JcEL6eRK-1X\0f,86gK,/UP4f+[dP=06K70RgG=f9M.LLXVGT
DLD-bd+TT.RG<K]PD<9>XG:TLV+d3FZA./\/SK^H<cYZOT^>D;ZICd+X107X7ab;
.5beZ3Z9QAf?^1(-3L@KS1<Z?.Cag<?&]-A[fOB/46e2:eJEB7_5=BL(BPcEO,5<
VNaPVKQFL\8]IHf&JY8)&3B,dfF]:2BJcH5ZHSP#SW7g@@N<S4P3B6Z0_a<<4,_Q
1XQ6A_L10TO80gA[[N,/EM^43VdfUGBde&bWH7U<5FJT\8]#EJW,YLCP63gU<H/a
VD5LP)C+La_+6^F9BA^4?QOg+7?NT55<B3(THEJ+;DG7g&6N=<G\6P@^2^f].4HI
D9K_>B8]gHfSObD:<b9K5]K4.UAV_S3[6EOe;(>)^UKPUaSASIV-)\Yd<#>5LPY#
[T>(^f^Kgg9e7bS#R2cA]XPc(TL1K)O7McOSQ;-->-M;,^P:aF36SJG>^^/&UOe=
c/PHUC-eO]3_\5]_f)1>FCS]aP&VA\K#CQT+/Q(gPI.@39D&ZdL_CEGCM;3(2eY&
&?^&K);6I4/E632].O]aZ]YV4HT6@I.\-;[/=PQ9(aZS^3OK]LER9CC/^fWa\fIQ
UCG[=cDCa]H57?,1Q/BM7J]TB>=<Fe/YLNF@;CE6@T]OTORATSNV+Vab->F&bN5?
e:f1:4e?dJMD2D>PK7.-CPA5T:T0&>S\K6P=CYXT<Ge-<2B&8<50/G+@5L=AG>0?
,)KOGeG&OD,@>FA>Xc#4fFJ[QRWf^TB?RYKcE^;gd(^O_R:R2ZKC8Hd\A).,:[.E
0Sf395Qc/gD1WJgd7&>V;,:_-A6AJQ\F>(?+cc<V6YI5bE.Q>HR]:F]_(;4M;P\B
Q][4[9-2^c<)VZ+3:\E:4WJ\#ZVO#fA)8HIUIe(\IbF,?ef6MYgP,YBg220Id=9I
[-E7O;eXY)g?5;\JMb(0,f4FOLY\A29(Sg)HW+F6-,)Z)eCb)>4W:&Rf3T74S_b,
ZV,c8f:9+c_d?/gg(]DI8<UG\BaFM7GXDaJ_BJ2J=UZFfP<22,#<X.ScKZ,c[B3W
U;-Gg#S23:W&[U/=A#MDSL,,6]e@7P?+&EQd.A\4=6H+cNH7UO1HRZ/H,Q&4I0-F
Sg0TRGGM.F>aZ:GZ4-RL:F)[2d9,-6^M;L[MK?=G^XW-M[U?-B[bG1Me9,EaFX>8
WL4)#MRJZ=)ES+EUL1)B-d(Pg.9AGc(S?fD,c>OT72]#4Z_.(3I31+X3(BH,L[J\
=]=b2E.VBUYGY/A/FaP2=+?_&:&JDR@ET?PU)&C=_.a>ZNMfcVC3f_,)X5RFZ:)g
@U8fMW(f=P>H2;RgQP4APXZA8UL+?P1fWTP-f-TVIQZ??e+FW?W;0>VP>/0YB##<
Hg0KGIOVWS=<VDd[>?8TUg1>JUGAJ_?e@BEM<WRU?D4ETaW=,N7gEQ&0fMX9L:?X
L]:F6AMPe,=eE#G-5;eUD3NPELUX2=K[gS[D:1JHGLZI3Q<4+=S,@@A^XT0HO3,6
gb#Ra:2QVb@cXW1RK(M>Ae,1P_Ie/VE7(_\.?2bLRR?<PAd<QbRC8A\TH>^FT/?T
P-Z)<M.PcW#Ra\,\39YfRa&H?/;Ag<6M3IgIL<XLQZK^ee^4>5[ZJba[>A(=F0+C
#:57&FG_MZO=NQdDI\/IBZU1#b/Y+Aac]-NX8abc?36=A]f#XMgUI(/?2>_B49D9
IUGQAc-DQSCfYaH>ONgE.8BYb9&(gD]AS6D]V-??L6>cIgXQ=P.921Db4M>Z4E+&
_c.C,N:TYCbD^IXbV^.Ae=,_M[X#@@bO+1X-&&WC.F;KJ?7[d.Z;CLeD^E]X+&[7
^>1257M??fcb3,Ga2_RFTU^M#=-@A/F5V6J3B\(C?eZKLFgF8ZVHM.>\[g^AI#U^
EgTY,,dg]7@ZcI,Y801a5_BK]c+4(]@/I1<feFBFFA:>/.U6]1.cS?9Y<^QgL.QB
6^KccFH<[&(5<43fRN/2#OA)MaXG<C6@GQ\a;UaCGEdVf4,M-@P/KTA:/4#3fY>C
T/7YFKd(;&DP9_&;dWK^OHcP&7LR0cMH09#ZKgPQ;P(gB&D/@.<d;P&-.RONB:FJ
fNQWgVSLF2O-E)J9CX@CYMb<V0X-_fXT#\g_aZ]D9LHKWa)9,-5bQPUAXX9GQOP)
gHT.KDQJ43;Y:TZ1OG<#=8f10(5=,VED7[acgWg#\N,=P=S=&&CN6K>dNFMfR@8N
a\)V60ZV;g=Y@1ULE7RKVX65K=FP[KMY,/P.;BZOR?=T_)J]9d[+]31>>,K-V597
3_^e8?e@EGR_-754ZVfGY_S))^AAb<CU0<C=;3?F11FK0ETS/0D;LFY]DTIVd^#V
(4fQH&C^\@A>\<T[GaOXO3KZOILcb]3d@59N:Ae;7G2^Y+<.R,GUIG[;eN\#f?&9
;bZD)5L2gb?DfT^1d0O1-\ddO[ALf].([2[Q4Z;]Fa[(4&2(E0_cOK#Uf.&Q9HLM
I;0DPG][.#.PC(I5=H_2=^+]A],DY</V2,G;1HRF)NI8TCa@S;c>]\DaIOX7XaeV
74WUe:KQ\E:g]PAf-KW;P<I_)^X>0SOP:>:aBefX<f,fJW))Z#.OXX>1I2JQec>W
>1gf:e#-QQOVFLU74((ML8.bBTUQI8R.-D&g([@/PMCN[.I:2I>A.CTMHTIB7>>e
P-KYM]^SBb1eZ,Q?dJ7g&W_[H?Y2S.d)@T6U<=);5^g52((V@cN[bFd]IAPN<XAG
NRU35<M/a=(c42;V0EY@:1O[1#>cA-UM.Ocg,gKgRW+:F4_)G:TG3]35W@6BW;R]
2L1F3M/R@eKTT=QL6M0;WK@[_SUV8)Y@]E9=ee5T6(=IX-+=8:?_S7WL(G:1;Q[/
AAR[>e[XYV;L^bb7aJ<8-(Le0e2YaOKW=GV<R#[_cd#IP157/9IVQb70\LfIA2#+
,Ya^^?Z3IB\>^,6P.5NO,(#:0@;Q/P1WT&TbdGV3=b84Z,BA5ZcZ3?YbR2:;<J2J
IZc#P63I<[&P3X5GU:2AQ_)\3SdR3QX#Ed,@],(I5>f0^g5W<8?=,3C^7I<6-O.5
JD;UCSHDN0E=:bdFb)26Y-_XP19U@P(]ZY[HNE4d6A-PgHfW+Yc6Z_I+7H0b9,Oe
-_&&2IYV2@FA[-6-K_,?,)E4>4dKf2[CGI41T\94,I>d:ESYGVG7[.2SA/?gL4M,
W09JQE7/FfFGI:=2B_;O[&X@Q0S;J7O)_Af\6J89V8O;P^+V1gfOKH=J];)U#Y@9
;W61/(RP)5dB_@/12Y>>SAFO@N?3NQ5)(;5DBL:<SCeZ&A#P>BWS8#];]MOdDN=6
dNe0AWgP-fBF1&+KPBV=#RF(<XQTF#B8-8YbAW1M<8:B[dgfOV1.)aL;D_L&WOT_
<7BOG36NHFW3c3T00K8XaaPgE=d.QbIXX]9BAH9W1=]VDYbZRV-D@5K6IX/fPLI?
L5R]4HONB^;QGXB(7S\KdA;)+4X@C5A3XACY9g@+Q?>b)CYD4_FRZ#PgaG&VY<d9
=UJQfX/M<gZ-dfYS-[,Iec/:B9115XIe509bY>G#ec8.8MP]<[Q]IT1VEJ-R20H(
N>@ZUg.5/(a[WccB7a26TAHacSdXN^V+J:\HLY2g#:,24R:(1OSM>dEVA:XMfZD.
O+G\baQ/]&1G+]Z>@989KT,X8R-93(=1>L-#?TP:)V5LQ62G#N5H#^PWYG9W>VR@
TMR;&L-(9JYGQU>3VG2S6Bf=]@5IH:I.4+#EG<C,P)5fEWONN<&N3E8?9X(=+1]a
OXWFK<ZZ;.4MVM/0W8X7##cWXME0cUKS]Y/G5^,+/AZLQ^c)R\b4g#CZ&SVA/EER
0;(cQeD#6<1_Fg#CGaC.g2&4,DOGO/P@?LbVQDE+H\UUM66(_C#/,W2Z7CX);N:+
\-5?,)XYJF7cNAE(PP;>^PD9+:F;RO>dJV-@HV>#bLQgB#V]?#QB(De+4@OKK[#e
#C?V)+2[8DgDCD:g<7SdD1.HG\^+VG=2Z#LMI.R(NeM4D(GZUJJBB7Y\,Ha/8eAE
0X9L<a:49Y)+CI>K@Xf70);d99AFJ/7\6Vb.dO_B1/5_;T[?Q-12daQe6_F&gKcV
_gS)X(2]ZW3?F-=dVLVR3=1e3?.@F]3O,M8Fd,5dBdF5#<5[X+44],67TJW3LQ@Y
)K7TgcK.W#QD]6;>&gN]Y.?EH_+/?)WP^cKPT+Q.WJ5A5QE_7Q.0OAK67^13#Z:+
4_=+0Y,YEV)BS9;=R#3=?K(83LSY=TM,UHZ;\Gg5VNbXa==7FJZOX?D,BA0g03@+
b(4aU-LTM2\1MHR5#b0E5-G(&VOVGQ^g4BSb2]PBROfaP9L?U0ZLaf.ZGSbWbWD[
eaXN?8?=Fd1KP@OSU\Ye<TQ^e^9D/]_.4).,:<796WT0OgM)\G4.a@:8#XJHR&-K
EXe=D#->>_GEF0O:c5RZU,C,SU,\bF\Tc6bHbF4[Q<HfXd;;_c81>[#8Z(I859G#
.\<X=P;S]-+SBBK72bI0eU.YeC3L#a;^(3XO8b6^]Q&Db,.g0L0GgZKIRe7\>e/N
DI8dI25@]815Q)<#>BN<.]_W/70/-C7N[eT.Gf5U)gIg/KYGA25Z>PX5;4AA_0;T
)5>e\X.JLPWMGRK-LR8Y?Y-E)T7YHN/eXbJ/dd2Y@)7)V0-WU]QT,SJfTA#c#3#\
[_NcMOB:ada(K4Se?UJ4[DM8I@AACeWfeJ<;N\)6P?/GLKEVb_,ODE28#OWJ=Z<O
Sd]:,d-[K,UdAT>_D+N_MQ(;d5S\LD)=;__4-<baC(f&/T;J_a:#_=&b/ceFg3f)
Ua^LGg&W&bVc[MAWE8O/;F/LRG>G8=P8bPM+7^^b([#@gBG[H,0]b2DS^#Z3N6Z1
(V=A3A/Y5L/7K^4VCeTb4FV(@H/E80N&.Nf6OIVWG&Q>G(UN:<5P-0SfG(3Jf72V
&P;#-Q)QZT)1EX:D?WGG:=::A&/[<2+[>&QKe,+-W+8_?BZ8K<36<<CFVI/?@K/7
JQWcb&[Ad4Q(CHPa=6#43aLHW(H-]fFNfHcQ,\?\AgXQB7G+[K^Jb_gED(AA]A.4
+=&,-E])U064D>PVU:=7I1IO3AO3cHK3^I=:EA8[_7VX8-MPDF+FLcdWf]ROP[I1
_^7P[Bb#KENA&U]?QPMD\MfbUc^.,@IU3D1Y@BD>BaPZ^&I<\@6(_9.OgDN3^>>C
ea+>dCb+61e@U.-eI=P:TS>7#4Be)WY.RJ[Y36\/I/)TG@@R13Z3>(#M5CTCE:)a
D&3MP1X1)NaVS#?Y@S^TPgOd<Z28&\9+2&a7[8;TCRb6.(Q9#V):BY,Z)7&fM0/?
;bGG3Va31)_,@C6)S.=#/(1);:Pf4c_+<VUYbgBcV_ESN47Q(V<;C3^M(a3MBH.A
cZcU+TRBM@OeCKZ6FSULV47<LY@Y[/JMD+@3\P68\Cc\A6BGIRN?T.30QO&c:7V.
,T57N;;=T.U#?W,@bHB&3AR=SL,^\<]-4[X9EgPd:MFF7=A:;]C1TaQ_c#2fe\;-
2P/P159O=4aFAXg=-g#MXF5@9ZdY9GJDBQQ2UJZ:N1HU&?e<1\+GVDPK)]bBAX.a
8XJ[Z;d2]-HS/5;<cT)5\0<=2>f8/0>bVBA8L4+83_VO=J2=;c[+QA:TVe580e^?
/;;I/a@:SE&Q[M[8fLN7ZeeQGDFVSN[B\BYF>>JRKKF8G<a6(VOd=EfK/Jd)(0YN
+L,HHfL;U30:85C4@PE4.XAd()ZLO/I7g<K/?]\ADB81C+RbWAIVZBHX?e\3?TZ6
O]>DIbPg+dLJGHS>,M,6I?,D@e>HWPS:0&R]QZ694A64LS76^g/7SSd]J01aO7TS
DbXTZAeQ6,5LL90@IB262BL+@T55P2I@KHM(B1Z=A)R)a/=aNU0GGT^6gaHR=F6X
HE/LKXP_2U(8OX\eNLd>O;,?@A-ZW5GbGSKC>c-]gQ;;ObOKXT^IQNTX@@=25ND]
dYf==d\g<4)8+S6AFS<We)5@PJAO;4@cYWUSOD5KI5f#\7)N6f+gCdb(Z9+>9U_@
.\0Ea#,0OJ@FZ5#^/FfZ?6TA<W_X:(XBE(dbXDEeN\X4.9ZJRH+3G0.9f-SWPM_1
MYEe0b;_J7SCAIJL)I@.5SLbBIaCD>CAA5M0[7BG;8=J.:Z:RVTVO(7-3^78THM]
T^JFKL;_\1Y044R>H4V7/75S(:]DF)_Z06V<BC1c4.Y8d;82bU3[&U0c/6K-D76N
J#[\UGYKLI+P<)\ZP2AMISNT1dY4#]::V.-KBEFA/D4d+^:.fY\9&A[,DLW0/=&L
RTW1S=7+<F>2@P?EO]@DCENE<;fVEYI8R0\Z?+Fd8^F=2S[XSF<7E.:FFV0fg^14
HP<2^PC=PL#J52>[#^>K(6V,TFZa,Y<:;4LRdTD.d:5ZGf4&4\^WUTP;2#af:e7&
]357._[OR=E\9Zaf<)Q8NS=ML[]Y^3Ce0+,c].=1EgMebKCZ]N5<TTX(]eJ?UQY\
52GZVJ=J-W#ce41QI>;c\42aTI-[XB\FLS_B:=Q_d=H9A9&5)b/6aU14OIMOE2Ya
1DKfX7&eH[bLN7=XbEBV6)V0GOc\=+MMA5;g7&6MS#Ma?B]&<aRZ:[<>-&E8[a2-
)]aY]eO7f4aT2_#CUe=D.V6C.a.d_2)DA^eeMJ1-;_(4DLA:3ZIXR9HHVKSOc2d3
,R\EO_3ND70bV:@OH<_^d5DYI91[cNJ6R^KGR&6cM;c]Gc#=NXQHR.&^)[9D(9+c
>LDa#6@Hd3VQGSD^SH,b;V4(+&6:b+^JT?f>,,Z[G&:42^Jb/A,MCL(-R-UgIQaC
BUA48Af3EUc/:2IPB=-TCfg=WVIYL[#d42IXW,g)D)3J(AJK#\.TE?]RR?7f&N)/
(6dN6RaSUcD>G@9-YTIgF5<gNLg:9\d79M&:EK.Re.Wa)QE\M?-,abVb<JOc^I)@
W(<9cbYO8/1]@?cTR&&JZEB5]R-.G#&B.(^[6)7S<H#V4^\RMBHK;9Ka]>&S=09\
8LgCO<WT=FB5TYL135J<M:9MPbHbYI]Dc:]-[11@d_GAU^[13+P#\A&F@aNHPI&^
0IW^J^UeJC,]g^<?1O;?Hg57S(&C&YS=-Qb>.HQ>KE[I^,P4AWbBJ#ZaWTc=D3B)
K_MH2WFJTA8;<\86;Y7143W>S#18@V/U<3-QSUDY94\Ke8?Y9b/V?0fN6,42XJ1a
XgRNT)edJ[/4T4X&26-Wa3C^13OAJJG5c[P<18b7g[.^,#bH@eY(-CR8BQU,TT2c
^g^2_&^Nc7MP7V]?R[(-.5^W[T-EB\Bb4UdW#BfVT9+IAGR^MC#L)SGRY2<343]O
QAK1BQagN8_^\VSBYR;d82=<a;N^0/gd5=gI(?gOH4ND2:A\I?GY/?8>AU^9FM.N
:5@/e=P(.,D16^0#@[8;F?QR]5,D[6bL6JCOb-A,=YKOOfP\T(eU6DgF7K[4=C3+
Sc_RZS5)D2]A8MEQZG.1e+fN@\a##<b5W3>G/&OVfRI:BL))@.=WKfOCD#4:+-7>
^,0,042Y]C)HRC4b\5UN<1:+4C43CgYUAJIg(K)1KIBc8PU^1_ECQXKcOd4Ld@+;
a3Uf3T;\TF[<DO=#8ODH,a\]#O<\[deP)2-N7fV6RZ3CV3e-A7AdEIZ(62BbXLA]
^A[PJ0UJF5H4,=J>O<V-;69,T#YcJ<[W^@^AX1EcICe.DdUAdR(C+_1W6\F0WIKW
1#+ebFD>JH8KW;@bcWNCQ3(JWQ(J>fNNZ/K3[>EF=)50;@^eXS^Bb=E<BR\Z).:2
PGDC:C1L<0f4M=9IfE>/?3BX\Q<15[T26Y=BHGgK?T,CaEEW[ZX[#^KRT7GXM,=M
P6TL<X#W;E37VffbVYI&JO#dC,,,NRe0ZC]E)@)L=.8.;E7P7F:Fd[+M>c.)_?+3
A<6JIbJJ]WEVaJPY1DdXYcJYV\G,KL)QZ/Z8gN,<^,/3(?,eUQYN:9DbD[FEVfJ2
ZQ_\Fa[/bL6URZg<WEK^]YI1^:3+8c9\&BfGA8Z:^bS,S#F=S@MR49WS)If[35gM
[1XQgHMQX3#EYO-2Y#I#@.gM;Z1()G1JP475I8A5EV.@&8:N@199Kd0>H\?PQb-9
,#=[g>7E_bAF2LLOA;8MX)D<Tg>BXQAMfD;]V84Z8)371-:5UQ44O6H#=SK:;//G
VIbc&SBD_<A.BPa.\E2GC/=]/S8.ERQ:-HD2&],bPPYQ,dc/L&S-(QEP/]-^3U4J
IEM6e]YbWYDS@&L6_(da)4Z[2RYTL?Tb]D#@<()4[dDXY.0GW=@6^<F@=8PeZebS
^DcdX<PeK26JXK676PI.HQFE_9+CdC,M6Qg7I_<\WRUV_g&a[,HBFU6]NVI-8;CD
:J8<2Z_E/HJa91?JRZRF.HJWPRRR-+C7G.J.7HbH5(#FJbB>(?/]3K8Y,RRHH;Ca
=f(NdG/GA7\CKO1\IPGV(P0\6:)ZDX1bT[(d>YDGZ2M.^:/8([:aW):OOO:Zg.@T
YL&>bC?HO_JUQ[Qa,G=6-Q#W/;Z9K&HDTZ2cD2WTNJ;-=@J3fRY?]V7aKFA1R5eJ
^;QH3BKA/3.I].C8X>aCAFEfR=7E\Wc>GYYD>;T9-0WIBKfIRI/8X5aeV&Z_?LY\
^:[a6L(Rf@@L8BA#@b((>R20cEJ:XE\X=)>.#)a26]XD2;Pg(JLG5J<,53YVN3GR
L1Ub3&:B>AE;_:(Jb)dd>T8Jg1,M5K4F]:8_:J5V5U8]V,EB<?Xf@<VcI<.&#cB,
5A<FXK&9.](1\Ug33UWH-YT#-G^^N=Q);T)MIFOHP18b;YQF]J_?(3IZ.V1g7dHB
Z+][#=WMMGaLHTM;H/\CK_I0BJ-)EH0F8<a>MAQJ>[e?[2:ORK0aQ;5g/a2(#TK_
#ZKES.MgRNaF=N&5&F6fY,V\(X-9#0C;X9U.b2cX14FPGVO;&9W,.\/SQ)Wd-L5E
.f#AX\+RPK(H=3Y\78J-Ia\XL<b;+0]XUb]NAg&)5+=Y[[T8\D7R^-S]De03(X^a
GI/94@G--XYQ6Y8:T1<R?ZA3gc8?)0+++^S3VXA5-\X&C(J)?=<3IOg[=I)X@?C<
80+[(/CITTK9?HIe+V@6N0K4+WIO;_;D]c?U;1Hf3)=K]IdG2&44._aD:d]Q93]V
JNQXM6M[e7GeJLd-BM_[e8[\7^S4-^_ZH&0>EaS5FOFF9QgX&4V+_bK)E8@@E/\E
+I<+-[D04VI_[ZMWQf7G,#^9@21@fIAR6VeIcf:_PYKNQI:(AB5&1T7A7VIOddfI
LM>CbM7fHg[K5O[06X7#??)/[N+,OW4OBA<_0X:-X_S)H8F.)8,H(SG<B)@WK+ST
7C0+_GT:LI-ZOcc??().d:?.2K[S.;^g=3\)LL;G&\Td,MEVd2?,[gN)\4#>T3P/
3De8^X^S]X748KE+e4gFS^.a+Ia7PE#,:+YDF_CT3Q;;;d5TZ00SF3K0dA@VM0M1
:WD7^eAIGa4.L(cLgFU>7KZVB9+Ka18](_?bf=2NJH]:Z(9,?_A9g^?.XQN,\#H=
\d\Y,(e;C517O>U8KP=ZCZH.:U2O-U3TQ4C>8V&83CCbER:SX:>e8Y?>ZdMYcC6.
df0R,-K?A94[W/I;XU.S_W-[&X=?4Od1=c;g>BGdQ&M+dBG2aMQdCLa[OS&E:gc=
WSC4];P,C8/6M,QQ30#W+]WI8&C<Q:[HYRHgPO15Z&&bJ(I\W\F7ecH4+?Z8<Fd0
-#AQCF:We>5[M(FACBL64_#6X@\IBD4d41/^MTQGaL@F#P5.9gb3)6HHPP2C#L+D
e^/Z]U>eF.;AD0(AV^&1IS@P_aZ_:fc21f1_<^dBVD8\9PBPUb9F?+b>P1[2(OA&
D5M(C_4/V5Qd10(f(\,Y1KX<.-7J0gUD1?#e=&DF.Z8-@eUZ7O/DK:S#g8NS^Oe4
TfG=&8\d5_^0f=0],S(4AM3Q9HIH7YEF:6AJ+;?Dc07I;X1aQAH5e?Q5\9PODcO7
dcNb-8QJ;_e/BK7DK733YN1c_d[=BPD-1Vf:O,de72.??IMYH;PU+ANC_S_4JI]T
&9HgR+C7>,UG64)6c[_IfeKd-ZRFYOa(URX9+/dBEB7c\(5O^GbF47SW(LC82-/Y
45]HBbMMVI@6IBMVcOSbS-,O:G]6C28f3D;VN_1O0ICO3#NSM^O97S:e5cY\@#3e
-L<\LS:[Bf)E@5VAMSEBSfd5-X4KX5Wg6XAJ;B[I@:]D1S>^/><1\<?;7eO58^9b
&J49;TBRP:A=3W[KN=_fNSAK8fXC8J-<##1B#24X5T&a:H#</^=PfJ52T7#c]QCQ
.,89;89DD<=[62JQ:Ce+PRG@Qe<14(V1@+ZH_aJTP1>+T]3+X/:L:@CE3]1)-M26
/<2P[.G5)4NcZ8.RP][R/+C\I=1VX1gXQ:RE+35L]0@.VdAMFGT;NZB(fCPe_CZN
XMX@/I:>4ATK])-EY0+Qaee<F0@7-(ATLM,CZ>DZZUWCd&;gXSKE+,SAV?3@XID:
L?B_dR8:SI\eRN2A=bL&I0(A8L_F5aYQ00=;e8-YWE<Lb&ReXSP-]GO;dH[XHT7_
J0+=f7@c<g23=g,Yg283aZ<f/9F+6XC:L530HOT&\cJAH4f.1M4]77&3W6F1G]+>
/EQ=EJC7PL((L/N#5FdSW;R)eOI(d0c.J.M.=9,,XZ9,35#+BMX>]a_9g025>4De
0X)PVH-G^S8D?VH#KV)<_T5UZ?@0=ZRX_CSg>#Z/CK<D339@]D+H89A))S_N-Y4[
P&0Ja^O^&6U)MN#9)@fGDCXQ;8dSM:\YS)F6Ig_,ORVLEVKHZKI9b[Rb]^8;ICW6
8fHLW+QY@3.)aFX=.5e/6S&VVIO#-^b[E]K>QXT^&[>4gL<c+0ee)Q\#VUF-.D?L
3_X+SZ11?HCeRY=:YZY>aN3eH]ER3A+?<9&]W<,A80c2YY5LT3IUT::HYaQ-EEI)
S]@1#G_Z9]=aEWSO3gLf:NRWY3_>d0?aR&]H[G0A;b@57>NL-?276FHY6;^[XSDb
-\NU9\f@2UU(3]P9AK>dg&TcSc@ebF5VIV8;)D)<gUHERC4(G:VX:?VXF=)]21b.
>IDCXPE3^d:BF#dK0P-c@JH\K<U7b\]/./J3_S[@M?15Y\b8-+RJXFe^=8ac6;]F
RFUJTa5T7:B:B-43\2SLQ09+;3;5VG(AGS8BE&ARA^7>#?bHK5d(.PM^eK@N5)^V
a/B(PV3^+d@>H#YfSL9Y[WXM:8CP0)RB/FSH1B)8QLGd;)UR+Nb+CJeP6G\?b(G=
(&@=.0:,fO9+]PO/G91<.<6+UdTH)gSX:-9CTN2G;L)M5gJHJV99JD^Oe52M@6-U
/6<NQVOTH<U)9QC(&9)US8O.QaL7W^C1O/4V,?;RZ0O<V/,LVZEJ&-)Z<+e_c-a:
fFN1[CKR2)]4.Q[SSD3B&_(1TYQaAJAEXCVN49YT:OOJ0J\EL&M29bP<4YgH+11g
6Fb(,#gAHU6dT&.Ef78--ZH_7+;S5H.V\T8M^-QU@X?\XCaEAU_8R1S_C?IQfUN#
9U5:[:38bXaI,D^_>E+J64JGd7>SP/]9g]HH\T6?c9AO;QcDI_MAe&84Wg4,;T33
7/QDX1@D3I=gNb/[Yg<bL72H@W3[8L@4[(,YWPce=4SH.TD]EA6<D?._3Fe[)D39
&8?<Ke90b,HcP:UP/PgI)#K,?FNU)O+X1caD?+SD+]Q9Sbd^WRcGQ)7K\SeKb^gE
fQRfEYOEd<,LTVIM(_dU37H6^=baHDA]PF(Q9=Ag[@g5XMf/W,VM<:Z=6YGWBEP4
a1d@/_QYO12HHZee\.[@2&fEHcNMJOdg=4=&^e78._<a_P69)866Xd\^?^J2(6Q-
R+-QQB]RG4AMBf?]Z9?AdUf8E:EM>6=a/TaF6OD5AOY,eaf3OT8MdcU3N_W4ZW5/
Q@R(P)1EbR1@f]BY,Zd\PL+aO,W9bg]/P73:JX&0/e@J9^VUT)\LT,\&Y)Q5.0X0
:FaHe3,YHHDabC3#NQ#O5C7?JTCDaXB,330fe,Ve(CcYHU.87O33;^8TY+K9G5e3
89dY+OQKPP1eG#O5Q>^0fP5,8c9?4VNNKg).PeY\bQBWZ2,W+0;DVafH(D:cG=Q7
d\Ad9&bga?J>KYd\K2@9&LCI)M/Q5)6ZB8QgYR,eLg\cTG-LX?eTd&K:bAG^gX3<
BG(fQgXMdDf_W]D/3#CW4R,]U5@6J_1LQc_W#<f]NUgS(?<#MfCT<65?FD;55AdD
(AZ/6e(=ge(OYEg?,B+#/EU/)=?X0JJ7++Q@(NDaV#J2>.\&U(3NVM27<dgN3Q;]
+/<].aa+^KC]WFY[ESZLYRI]4C27VV1b\5MQ-TI>+6^ZJ8>MeFcMc&KHNJFb-YXU
@:5Hf\C:OG>>SC9F2UbEfg5^::[N)g8J.Zb-\<VTd9__K_U)#0.Da[A>_7E=S8Q6
BTcU5#2UJLM]JS&A7c8+dQ;S?,0[^c2<,8^9L=B=ePLWFe/^I[NBNPA-Z/?_,L:V
fM\b1GA7c[,JbdN2,=B6[@C9[C3.(7(8Kc^FZKQdb8D5He;1YK6H.9dZGB.COd>M
fE55(<6g=39)Ag@8D&B?b[NR3[0X?_b\CF02S\e_8P(R;09I4?4E0>9+-&<CbU>5
MgdL_985W\aQ7NR7dTc,?GVF-0?c;A:4g1.Va:Lc(Lae+A91=f^66:NR7d).eQVD
1/.V8UVG;b&)Mgd4HD9FH?eU)[(g&9bR\A>.XR9_e8Hgcg0A^<)7.WNK)V]C\#H&
a5=IQTOL0UKX[]06M>=eM?VgJ7/4?_X)2.JPM5+I0+TR)S([:+X^02?Pbcd,VO1X
a]f/M3d#?Q1S-FLL?49?eVQ.[@<35;CXG0c+5KZ\#X091eeG0PY<;NPbJM1S;caL
\75bGSTB4MNO^cIT:=Q#;2)GI_#K[AV&?Q>JO@_=dF?OF+BF7Wg(#Q964J-aeUD_
AV_CPI;?^Y1C6BE@6:UT\,.1<5B,K@JED0N/87(c0-5>.3F<+#Z_Fa5e#BBbdZKZ
ON6cHXP7IPZ[EL08LWOFEWX2&)BJD3K]LN:6E<;2KJ;4PO@.J8TdRT];2]W7EHg:
O2TH(.R2]D:c(R2W-\I#=E6<(@ZRbW1fP_3c37EZDOG;BDOFTBH#g.AE6bD>7b2V
;3.:77[WO=;.\^#;ZBd0HJ-&6QI:]a:K8E(4N,GNB1Wf\7JCKE?K)(NME.I\AA04
-@^[2eAB?8BF/fY_[Q9#<bSK;.5OL:9d/.W&dA;;]H+9/bM/04J+1.UAg/_?da=5
EW8d@BVggP(6R^M=IV-ATX<)VP5\36aN,/E1W5bYRQ^62--=(&I/FP4aDE/][QFQ
0eC[4YY0IE9;^O^L6dX>GdOD4_7cUR[0a@7K1YC=[-gb:CK?8FJ6BZI:MGS6(S7?
E9:/SOE(6BXTYV,QU=X2K[?S).;(E->U3XOXA41C,P.=RC_NUH<;eX_9(<[NJ0S?
fC<>9RbG:[PF^VOUX0#a-e-&PYI8(#T/4DHMOKLL+J.S4SAAUfJ=4;@C9aCbd;BV
7>)a&a3H@M>_A-EQRfM8/C6P0CCa]ZVE\EaDUEO,ZJXT].OUGW:^ceH7I(E;/c6d
?0>B/W>(XF4RT7#;AX5dHI4GI]bg=0U;&cbP9bGaR&b#6;(P:K(&WJegF101R]08
c.L6<gW[51X#L&&<>A,&UE09VAH@/adcUCNGDBCQC9MW^a#69\M@Y1b]:H+@[c6A
K.J384,)P(H@BY(ed</NISRV@7V,Q>MMaY1BI2YP^6;W#S,E;/F\IDWF<JR9B>g)
[2OC9aRe2J5DIbS/8]=U:W0_Ng1g<?YH/gVP5a5a:6bg+,9LW\&^;#72U3FC-VW-
O<b&(FWf3L6;gS^<OG+251_5W[40C5?-M9#E7VHg,P<Z55MJ>ee?>TODNSDd[=gB
Ded5K-Hc\0;d+/.ZB49)2ENI=4X._Nf_/G\6R^/(>YD9O-A,T<]?UM718BK^O)JT
Mb[d==SYZX]IR3J&V6gLHQ?c[\-=^YLdWZA7a)UaCAN?9f:YdL=PS>BNPa07<&e\
Y<B)(+C&]6G=A0G972\bB[_0-^a8)4^#I9HOIG:>eB<Uc>9dK1a<;;6Fc1T2\]6#
]<S1<PgK+-YAKBB)+;Vc=?TgZ91MC.B?50J0U1W[@##M3VD5f.6HU,0H?<6@&E\N
_dWJ(XIM<_ESE6&[YD4W2T_K-TVdLE^f^D(]_XFa]5X0Ue>],\F9ZVENV2U?870?
+/1TaYa/C/+,dHGE=86b5&CgW\@3-3d@QMG^Vc\9aCgB62M7H0RYJF8<_S9H\WWc
_;1F\.E]I36N3L2B2bAGf95g=)>d_cZ#V_FQPgDa0:E.S>+Vf5ACg#;RfL1JbL^^
(f:O[e;LS+0TfX>c@^5=C57B&M8VD6RLg;QgVdCQaNBXY^DW4c5IN@XV<1I5ee?[
?QafKC?VKHRN4V1.4A6d1_gHg9eebS.C5HPaBK0[Q@V4eYG-]Y8X2)V..(>XFH&b
e4J;T4M80YHQ8<,YAGY0S2_eX3e_^eQIB=AO(S]>+MZFO>&OVdMBgLQeXANGeKQ2
3&WeO=G@(Y:MWPKg,HR(TLC(PeARLE9S6^I29?G0QLGWI-0.f9JdX>-P9b-1\([.
6EI-IDJ)TAcbOeXQ]a;<]UC()=B1;JZPQ7L.?M?_Vg6GRMcSK]PNK6)dX&;:KLd/
UB<9TZ0gJ5GbASD\]=BUI.2LDW+^JS&<f/A]9Q8:Y-8<T/M2EH0,.F]20)JA0de]
_,PY<]ML8FPd#?a]T+1Z)_aZ49cf3[W&E2SFP#P=(DXV=H3>/<HS.DC5LMPSV:eN
-[8<G>@>70^?;Mb>@64O.(US=NHR)>M_gJU&M3+]3(P8Of>].Ac2Tb?=W.DRXBLF
1;4#V(#c]W_QaIWLa?K2:AI3fLIK9Ff/g^(CAR[+OBNG<6R[>#Wd3Ee^VQ6Qc.[4
,B0R3LPE\EcD-+S8Y82I6;d+\YS19ZD>ZLNPBOJ)ZZBOT_V0B:S&49=fHM_A#ZSb
3L79Pcf^_D#QR;STf/O8&CU_97#3HXaLU-D4\7BNBTaCY_##NOCC(PQ>,2QYC\(g
G.RRQAB#YXB,?Z+_M)4K([IRHf]ZIVRG_C,\@_]RMg[X[B;deA@7Cb^)f8(3P#);
c?8F\O,PA,If&5XV<H_AWT4FP?8He\Ye3EWb8U)Yc2fS(V3J2:BVIg^DY[Le+bbC
Fe:E;HIG&(=B<(9KU6[/agO]F6HY&R+E(T3>[b.#GT3]Sc=/Xc8,_-4Xc18GJ[FU
#)I6EM)I(>E^^6[c+:04^P[7WB@bBJ5PeJ,T(3LYXZJ?NQRH4W(ce:+G[Oa2DH[Y
]>R43@:.Z2>&>G_[RdJK7^?eF-2II8.QO+J:4NFMN#S=6:e#T;L_R/COVWNIeGST
+_PGTN_=+8+).\\[YI7b\O\D\7\1CEaB[A8HYMR+.PW8.:6WA@bSD#9,TY-7H?JP
;5056.DBFXT..J?#X<5;LI2H]5?fB<#D2#DUDdPHLMfV80C=:;PT:2_=03ba>9]]
fQ@ILH[U@;0:I>,,)85SF<OS@N79,Y)F@bT(I=K+PN-8.Q(44&1UEPd#X[HPB/S3
e9.1[KX=/NVL:(+Q4.B54(?8I]Q/)LN@ECcRMKC=XQ_O?WM4USAJ5_NFAP-TXX8T
RScSX)cE2E11ZgZ:-+a//2KV.=+e3H0Q9RFAE3#B<@a>^e_3Jd7RL^dZ(DJ<A@>7
0<WCaN3@V>M,G>dE+Lc.(P;>aaeE3FTQU_F-Z8FHV6/[0?M]K]J=@^/R,T)_U&+e
gIEZ#TcJg5.S<8H,UEg:&<LT6<QgJ]AK/=(_a.W-\L8WBde)\gEG&HF@fF@L:ZJM
-:9aHKGd6M+GU?\LDO>;I(d/Ac)CRN,75dbN6==EWY9-dB-#cK3><1N?X^PcW[=\
G3U1L4VJAF]/X(/b>]@X:2A7J=fPE6\QNC46;.7eXLDC1>,X.SQ(0Q;WgKL3Q0RZ
BGEa+AOZ7/+gaKgLFUKTEaXPGdde=+J]bYWAEd,MBE:A(CMHN)/Y?eF-Z@N?:AO(
-^WSW);,>4N2E(WfHe<@WG92^>;@SRO4bM31_1XJ.>Q^#gK-A6bS],eJ<74M\(@c
=Z8c[cP+,_,ZgcB>STMU=Q_bF)UO;4CQO2<>cOR@,.BUP>Ba&=1Z;=V2QJ<TWcR7
RKKg6c<I+T-)Se0FQ2#;NZbUQBg2))RS_O/,XJ[f6/0]W[SVSQI-aQGc<KH@B,Kc
#YIH>Z[S<2YJPbV34Ba7-MGTN2B,-(QM+C68&.9UbZ9_S2E(:R?QC_IL<U+V+/W+
UbS;G:_bY_<A;M)N5^bYGe@.7=0Ucgd^=GF0@UK,EWQ25UcIEbA<LRO#K:Q3W.64
D8UW;[GaT:HD@<>/5ePU:=b)0S>GJ(4Kc0dT:/C-.Pe7P6Y\P]<dZgY16(c^FECX
Zd4#[B^\9Bd<4>Q6JHBTWYC@7PE;]V^g2Kc-f([[T^L\M0.g(\c/561+WWT@C64^
Q1X&+OgE3R/UA_8QI<HgP+PPdR5fcNTCa0RHNSJ4.[1aUU][MCS<,I76eMY2HaU\
=W(K,f5<fJ4V8g_48&g@_2,-,7OZ?-.M\cL?+dFa#^FO8I&We,(>+)V]bK6&Ff<S
e^XU)IVe\[V4RI4,ADTWR;VK(dRdW^LED[gCU>dS8+]:8Q0O&&;dRZ<MBFEUOYP[
cfLER;CAcY+,CE81=<2TJ.@)DC4W3OdV[@\7)K;6Y^HT<:H6a^ZLFA@>BF@KU4fY
cF)eYAAb01Aba]L9-,&X5/fJ1)/V<aIQ&((OJ@^fBHcDWa:/]Q+0PJ-\[gQ,NdO7
=]D&URR^MV7<0G8/#^X4S89_4OLP)IW2^=K2+_5UH/7]TR]f/YfG]VMLb1MD-PVW
:PJ@QZ+3VX=K-^L8,X>/Z(HcA3;@G.[UL./1I72RA(5+8+f;WMSPD&dIA4?WTB<@
X\6R5_[&MGfC@\?<?ZRPJd6R5;ReHR-Of(>+/73S+N/=)>C@^O1U@IIN__#5c?XR
MA#G@WeKF#-_5FF1;1MgSL#8K??5EVNY-OgH2FeR_((;655[Y(-aKda@FeSLXUaF
>@>c&OCA/:-&^\K1f?3:/@1/b@4IVJ9gOK0M?442;O7\BeOY7=#1B;ON>NL]6:=Q
,MDC6.46Y1,1gXT/>&+0\=5;Pg#;#<J8[>0aJ\JM6gCPC1:NA3=0_8)b)9(JO&Ea
TDJHLX083WC=Le)GI3R;PfZ,PDJ(@?]#J,&3<MJ.P>J1G2];:03a)T;K4F07;fVD
S:bW>4A9+ga7]4g8ECJFC?cA8LR+PWB?Z3CUYcCQ3GN5TfIU<(<OfL=5&e[:^/,R
K=K3CK\N-:-U\91g]fW?60?gI6@L3VX3fgV928M1EQC#.03(5dR4,>;#GGI0Qg5e
]LI(55G^5LQTD8PgVMUH9:OQK+aUfJ92.V_S[;N57PO<A2e.H]c:,LXU7KB))PXX
48HAaIaMD5/d0APJIfGe-D5YFc3eWFU/3@[PFHIf_;K8UE7K=N_aNcTM+=+.LS.K
H98TO&fL#I=&-f;+C:^G_QcP&MW^3UADK2)d?e]c08Cd1-7J1P^,U[0/ae)d090c
B<47+f[.;.(?bW<6#FBA23g7[C:O&5@A./IKgCKG]9fO_VJ/#8e9?a=[EHO]FF#-
C1PQ^c74;@?,d4fCZ-7fBRbf(f#If->=2=\<2PeXJNb7VOMPE1VF9T,904VJWS&a
1Pg<Gc9R(E(].VTJ5_;dQE\CbEOcZXL6G>eg&V@&KD=PMHBabA,/OVZa+T3bO+.d
&T@X-B)X:f,T>J9E992]cg@^AG[f>XO;Q])3-]K=4OX@RaN?JZJT:>09:TVa)@Bb
#WD7WJYF;g-C.I6CgB-<b6/@&gNOIA[3^-4Xd^4R;]F/=KC_+KL?T;LVRDNT#2]f
<CWH+6e[\6.4gX36-8bYcD_2AX<C[PKIYaA9DNf?FJ.gc3DbLOe>\:NSe_@FSgP9
R/#N8(b[-Ia,If@.+f&GF(5C5:/T590;JGbMITN7?GNO0EP6f(JN:M&,[\]cD7;N
+<TJ?3^UAd)Ybf.^a4C\^E&//&7,b@V1FdK1+AY64N.;/U2Y;/W0cc+;(W86.MOQ
UK5JZ3?V8QQbc@]eZTabQeWAQ/4aF9Y]F,N4bU&&5]W\AMNA./3RM@EC/K6,g]f>
]e6Y0FN>#AON4Q3e-A:d;ROYaVCNP0A;7c[^ZUW=@,3Q)-d&==Ag+EMF;@@IB3;/
6^ZZCVdBKV1VWE9P(P4T3OcPO#S:S9d=W>Q9/+HF1PDXFF/TPf60T[49#4XCTQMF
Y<GC\c6f2]fVO1=DO/(e/O5g-Md_e5Dd2^,@f+@_7e9CC,4@K[I(99#-)X]?c@NF
3<-,JYKY9WN/\4gG.H[VEegWGfa(c0I1dQd)\ed9M<aL-;DN]A/5K#_1W?\NAJWV
B)BP<dV7?C@_IZF7ZW]T?8(;G-5/06O,63MZP+HeHP^07J\=Q5GBHO;4X:fYV_G[
WC;G49T01\J>AV8]2,<fJgD&?ZKBKCDAF3F(GOc9N5652]TH@/:,bYFLCaA@&7):
H0YJSM0AMVR21N_65>U2Ad_3GN8UR=7@?SYR6=]TE#_[/EAQEKFS0<b\[+]?)9b:
_Z5+Z4_IJc]TEWT.8;b\D&3.);.<7LKdRf7=31VCf^YY;Z?0T0J8J<e/RHOYfUK<
S[G+Qc0;2YF.AC0eT.f,]cBX+P,<gRLBK5_-RRWKA3TVYBH)X^VM8H3BN)<U(;<]
;c2WT7NY>HSJ([4=TaP&Rc+#4#R=HaN.(KD)Dc7cO_We;e-8IGeLScE4XGW+A#:J
cHf(]7+#P[.0U,R7K(e@\?PHgA2NT9S,@?=?FJ_eHDF\F?.Pf:_X];4Y2&ES2gTT
]C&5=MUJc3/,LC7)JeQ#U84Yd[0R?Ja.(Ld/FOECR8Ta:1Uc^K+f&&-8;Z_+7M5A
TP)fGX3cYI\5_7Jec+_Tc(1cSZG83O][/?aBT39]=CKF[M;Y2-7aXB5+SY?V9aaT
5g&U-&Z.C[?Y<0dJFgfVR/d+RN=@RT7OQgKB\^M6]d.A2HQceTHDVMc:;LJVMbE[
T-\K/EL+)PA[Fe:gL3G2H2(L^N,E.9:#?6S[T.P[VXJFG@;&().b9Vg?GM+:Mb:a
)/OE4[@Rb\1?2S+1g95=d\McO]gb4aOJY8[66RF/Q]EL@@cf]8@]7HARQ&O1&-?P
G9\eQ/O)V4403fe58<e2cRfTBAOL6RH:-QVTf=_XS<I,NMW^Wb6-ZCPGgT^K6)(E
R4N8+=G4+2-Wb#-XUC.;9R#L<]R5F3<O2DXZe);7a2G4.bf,]+dSRO0?5[B\].T9
:6Q@9<SZ:))CMM0VRad(cB6NH^0ZaFB3IYZ;D;7,LE&Y2DNbG^J1^8J>4E:4R/\@
8/:TdH:]O&;<[=#FN9d.RNOXgV:D>(^L71=2MY:G0;.L^]_8XU?g4Rbc-Zd4/Nd>
YV,OKAdg>?T6H4[B:P\g]-JBZS@MWc[@(AJ_Ve>QG\)<DdS=JGEKf>OU>V\.Gd3U
_//FZF=/GZGPEWEZOUR]>@-04.P.d:_C;-6_+8faT&_Z0VOPb4\VXXJaP&)<I6DQ
gY@I<2FFbWO5f+-3eeCKZgP6Mf8A^G;PV#OYWNGF4W<bH(1X-R7G=392?gf7We0B
7&#,..PaGI]cAa#@FQ[2e^9A>JL^0],-V.BJP47RM_U70?;eTegMQaP#)]VZ@C7T
T3MAX4=FSN9VP8?1\)Q/7>faI],DFY2[90MD+:AS^J.9U70[G__,PL=@S/[W]ACB
(T85&[C8&C#C3RPIH1Xg^9ZWN46be?6/R0#GfS_CCfc?>]C;IY6U,JLM?82HO.EG
5aI)7OLNAVC]&?gbI-.=PNQO_\QH4-_PKSeH^&2?HI.]4Q?C?b3<__B[[1P@T,7E
e(,V&@b&GTPH8Z@\>MX;Ld]C.;MHL9][V[UX,Q38ZJG<FT?I-Kc(UC^6@H4bY?/@
U,_c-1dZe4\QV<-E^V?Y_M.DS2#EQ[18.\,XdMWJCAfRTH<52Wd#X24>g^@?4G[d
FZ54P>J0ZgMe]fa)E0c9R)dNO?gK.43&N>0eA?7S^bM.g>d(7]f;[eN>5C-EbJfT
A\.=E3fM1<Q]4D2/+1>_D/E]F)YaMA.8EFJ[GF:^3Q)@_+cM51K1(;1_ZZZ76fJ#
>C,c?V)R2A>IPS82P<7MJXSER7G)UZ#VAA6-a2&a.fH<V9A?TCTW]=X,E,.#:f]Z
O]bQ#S3XPIg3I#f9;1e(W6[;0T=aBKf?;S/+E>.L\f8&UMFNR;T-[B+7b^CWU3d#
fJMD^3L5c[/dE0:CbYK)Q,YX@64;54DSXS)E^J?;2>.;\d?A#-&U0GX<P#HHGUV;
J.(09F,VQZCDaF(WLAf5C::\DYVKU^5<E/1@+;>9_-DYaQ+2&S<^_VK_KCR\fJ9]
J+Z,:_=\92.XD&-/_V1&L9[FB4Rd>Fab=?M-K\d?;0Y<dW@1W->G<;VH1Y/aV23d
>[N>G7Qf+6=<T5=1T:7;G6L]K3>Qe@=c4M.#Z,&QQ4L;Q8PL>>:Yc3ODA&U>K^DC
U9(6]DdcTdHC.\\0McOcL,:2Y?].EC1[FZCK++#C5-bQVVA#.cHZT\GU.VN&KT;?
:98W+#A-EY@4(Tcf@=CTZZBf;LWLNSTN57NB#2\>WJX4(\1:7#IS<IeWO)K/cJ1Q
N+@dP_[ZB?D.;_g/J>S,P?SR\A[J3#.>ZW,QUOM4&=LYP=geQ;g7-)?R?S<5;;D+
03S:GN3JBA:BeDXEf@N9[??<-MOG^2/(OJXRMY\1:c3GfKTD><SZfMGL6O#B3B:F
3bMMM90)5YPP1ga,OW]e3?L0@>>e[S)WV(^_3,gG<F&#)/E3acbA>,^Lc&3LE8f_
PNZO(?:>23b<+4OC/39G>ZVDTF<&.Hg]>8FcJOe8B&SVA)T(E;^+d[&]40QL4D\g
_eN-9.ZK3J[\9)GdAK:,F9Q0RY._?Wd:=,f^0b_bW.2cO_H]e()VH@M\0B+^)-US
)E[+_MTacK(BWH9+EQ#RcL]N#a9#<S)VYOQG/8C#L:O>Rdd.I-?I/S1b2Y6-S@/(
W5XV\85PMRWQ/9:YAI@]/I]SO\aD_R+E8(MAS/9Z7eHgZWEg),9TM5O:Y]_Hd&2H
a52B/QeTJJ7I]fc:4H,<T,C=dXKPDWQ/,];FBNf\Gb0G](IaXAG<1I7I2a8<;GHJ
88I[bDX&/H(QFAQ<;<#HGG;9(7NMKCA);VSIa+GAV@#T,8Q)K1egIE46Q64>4]]V
:,ERWH1IIeWYA.?dKJ]W<49=EJ<@)6;ZI_^J9b=M2fR#:+]SW8&5+eeV(Acb06V4
M0XC87]P\HEZ5GX/?&DHeIJ2X]+N6MU10d;f001B,F<ecW<TS4ECY^TTa#67VLK]
D7P9TP8656X:fAVC1:9eXfce.S,EW)G-STLV:OXdQ7-M<daSW((X6EA:99M\-Q,)
L,f_OER#(ESD+XZc1Q456JgbafTaH8f=7.cZ&6X\3a-N2AHA2DS+L[;VPGIUcTT:
:/#D@bZ:(C9YT0U5JLRJP59FJNJ.([DeTXPDL82TJ2fA@Hd2IRB5#8M+>;F(^7dM
AgFT;U-Rc7+D=AHUO-OILI1></@_-^L-EKY.[MS?;d?/6D=fZI4^)IN+.H0.^Sba
J,O3H@S(aS5QY8X@4R]6(C8P8R:08)MF.T>2K&?V1#?<gC]J2^[27_\<J,4&&T>Z
7ZEAE=,[?KBB,F6WaS5<gF3>&.2dII),WB#JN[=/R6FM(9TR\-(:FK-L>QMQ/RO3
^b7WT,0O]3W4R4>b9D@XO4NL/M2Y+DX]WVE;D5YORZ,QTOJF[:-G:Z[GcKQ@P\K5
,&JaE@99)@Y-.?Vg/BRD[.P#3[Zf2fad]CRA_4>/.30f8L8-:+fZ,)NX8-E,XY.F
_K<4Z3CNgV0HIbObUaVc-?&=[S-+^OJ>]Q91]W;d4Ee\f7?RHIg3\dDPS;T9_c^)
N>&I-(=P2QVU9,bDAAS8X71/FD@^ERd[+E&RDTXU0.bXUJD^2IR;-5,BM&@NC;)R
J?G@g,=2.dK-[SEdH]=3LA=GfJFE1_#A6G2H+DRd2L/TL<YZPac-<;GZSZCZ);0H
eI4PGW^XC?R>KU<T513#AN2DVXRC#gEDZ==bVZ=E/S3/.WM>(O(TI-aV#g(WL-G#
B-0C+;=2FK8BdO85GWZ1\+,Fa/1>MP+E>8]?HN6]J@?1#)N51Q4/MQ)XS7_bGW+0
7--?JU3TX3BX3GP0T<^FYC0?b3LWNS8<b4P52e;_&JWW;U\31S]eHCJ0IX-NK/&,
g^ZgX9c@F]&EDHbRD;Q):YFP=3P)9O3IP4^\f;:PaSWK-6g#&>?58;N-+.0:G13L
LH\-KQH>Y8E@(caKDG1)DB,46CP3\XMC_TLKcg^?c;Y4]Fd9)HId7G@G1]\NDM9J
JTM+J[V[&KCPG=d4Ba1g]D&gcdGDM<g,b;F<A#2I;8;GFO]-5We/(7<1RW837?3.
Lf-O#@J5I-a=_>&&38BHU0/XCN_UV=F_ZMPD]&@FOPc6_1WSI;Zg2=]8BD.Y1A98
G.,E?&Y)7K5/7R]b+/3Zf[C[<T1HCE4@X]-[@QKEY1XR/K#@CC+[)JP6+Ygf3KB_
BU,,X93K4a:3J\.^MOga/ED:.>FEB/#GPYg)\GC=H?P?-__<WAR0AG[ME.>a3MB[
7Y>61c-/Z<b=f\2?W:3X3U@J(Z#\\&VI+cY(9NB0AEdCM&DZ<K-<Jd83TN=7XVG,
&-X<C)<-T.T,?VZZIN@gdR1TK8KDWTE-\#.GGddO[0R/,fW;VHIX39K>(1/UVI1)
DT9I(,e4&ZKb7P=1+&c.G9?]35d+M5CP?:dL?BPS+3]2&c;4N=2OX^-d1b@\Z2?a
&]>a(;g._KHM3(g,GX2POQ].1QgJZ0>@N&91A[U4Bd<R1ZO)a;B)#:-P]?()-8>>
@a:NCH.ba5N:O@McaVf6R]1H_IE;7G,BZ:SQ7J@UZbJ(3@+-1^2CE3Vc=^>PCX>+
==COe9K;E4NZH_+44B8CG0NW[O.K7M@+BCS)KHc?9dQUR)9ZfL7fF8//MRF0T5U,
bgS6>RS1ETcPPI=]abEWJg8W&5g>4>g?XL;[_.JbW+QUEF30(U2^C]?E2F_B6;G@
>CKZB@;1?6e)J1R;;EgJ.UGcJ?1bGUJ@fSCK,&1F8N/HeW:KgO^&g?.A\H7>c1.,
#?d7[I6]gHJfG2#X=M0?b:?KQ.3]-N<W]P@ggE3LX,^LAO@Z_>48YJ.P7NB#Qg8A
EYLERFdIB[8DD&+VK1E,UFUb0NR?Ve5DKFW+L:K4<F2JV]9_I;N909ZZOcHTOb73
cJB&TT/V6A0_ZT#SdXU91+K7@[N./^/=?dW60c[cf4RJ\Q.>&@3ag:#-TOGH=USX
<6EO\dA-70AQ?9fg2\?11a/\H+c_M7ge)J1Y4NHG.8SZ4QAd]B]KHQ:BWBf<.b^0
#P^c1;L]_fSK>,,?3;\P\=:O<#Z>OZTMTC7Fb5]FHK[c8@?g-MHG,D3A_3A:9MVb
M4F+\/OfN_GTG4+07@EQ1#RXO=\0a.(=NK/42]C/-C>&Q5?0CUKTX8]g,3S(Ca\R
&]Q)^;\<.[eNUL5E;:6=FaI<:IH?e)bOH&1]XGbFAOW^ST6-(13Z5LQ.\=1&,J>6
S).VHH9#;f.MgP8Z(FU;1D1B@N]2FPM2O#4/RLf<</[A4B,X[R^GY0R7D)S=)[a^
;BH1/(E\]Df?e[I6(?LIQN)81F-]Vd.OcM>/KA1@=V_8]VZf&FIHZLX3dP@[YJ:Z
+WB#JD33aI8O]0CD^7CT_BES@0PdI<:2Y-6d:I]9[>eTAE>?Z^DMXaS6PXRDV[8[
],D0ZaaUL\HT@F6,.6R-ITDWN&H31I8>7N-^J[MYC)0/aK\ZFb#-W-CT;<_OHE9^
.ENe2I7g3@W7(662.20Xa<)fPfY_+A^5XWV7]gZ>-<JcF5+TV4Z4A6Xf3SF_\VB7
]?CbJd#dI8)QOD[I;f<YcEd).PZ&7XCHZJ=74M-O+H=OeXI=J8LdH;\+b<.71Q2e
Y/bcTB\.1OO.<XZEeERP&LJR(Y?I(K;8QF@7b4=8-I<#6@L]D8d-:_J@eD>1>?=g
e\CO]_JH[/03ZU42]KW8.(XDaP5_/MfVM0bU>^7;L4+-[/R00?=@;Y[YZac3=SKV
IB^_VZN14MeP33N>S1bA?E&Zb&HDTc:T211g@-AK,CXAM>c#;R#Z)deHdMGY?gQa
]OMPO7L0Gc15H:01GH4.bQAgX@]?9f?X3.<__e>&54PEB?KBZf;a0)FDfACZGDA-
P@AX[7cPVWRE=cP#BWPUV,IYX=dG#@g2f(RJUF#K7,X(TKR:JMac=/26SV:[d>^X
Q#,b<CHFddERBA6BY_H(<.2Z;M:F+\dHG&[&95gF-=P)cF]cAX9O?HcgWAe+T^E8
&ZO-RB]K_@J(.Ga[-6#&O.b45<gMg)0Z/bFD;VLe6.6V2(\W&b]JE\2,b+MZRb?7
>9P6+DRP:64Aea&>Kd/1SBY7M0Q1;eRgbCc]H4g32);9/)QfO9P[?(a3N+XWf_b4
0]Jg00.b1<KXNgK,?W8[eL9,LY=#<=^gE\T5X3d35E3#gD/A(dReX:F-Q?HKc=]]
5WUK85Y@@Q.HEHDRWYU54/F[]I)D=7JgJ^,2Z?9gPXH#?7.e3a?RLVM@_N,LCER_
,IL0F\=A.0;U#BT[^ag7&&1YTdXJQLR,NC>g>>;>&+NZ5[)bHJ>4^d[BZOR?_X3T
0FN8ROW/f;gGB1>b]9@bD4EX.>H0b=a3Q#ZQ5S.PX5aM8\7PJ#19c[./2eeNEW5:
8F(2H&+fW6.^D/1@E6Lg\P[d:KLBOIB]1;,bWg]VH.I[6A3Z@#]AcT7VDdPeL7)\
>ZeZY<_@?eS[d?N-X&c-R_K&?)VI18a10XV62+FHLKb&(EBNS5)V_KZ7WQ;@XUK]
;e[3?^)W_bFfAH27gZ0FB\>U9=J(YZ<73cf^&S^NQQ-4fO.Pg,f1cW5M4[7]6]@H
6b]/WC5\d,;d0C[PW.aWTU8)>5;US5&]AEaQKQ]9&AgMKQ4?dK>6]WEU8^f]K8cL
;GUACX<-3f/Q_6\a2bAVR)5:V0/YY#.O;/b#N7?U?NZcM6eeda5\MSXB:d(9?=(0
Q/-38XZ:/LN;&I,SS]0X#U?;eFa+85XUO14\?gLT<[a+C;:R(/<12,6V>8#U]L\5
IR-M,DN]]8g?5=ED1AMW0AHB,#SOHc\VDCM@1=d-fE^b3_8Z05Mc8N&_)@;Ff,Se
,:(4Ec.6IHRX&b.I,ZIZ,OSD#:C]B7C(H<5-,#>;N@Hf1GOgP\0)b\?F2DB@aDR6
OA-d9[(<dRX@TIa.3]X_Q-3_KNHTOeJGE[FRY2_GB.\Q\e@>aeK[b<a9P^3W<Gb2
VAa&LC?YS^WbNT_4J@5D:M.JG=R@=QW<:776XH^6+fET9U5+V>&Z1+f@9>V]#W4N
,M524D>;].QH>E90T3FX6ET8cdHZFe(>c8a5)1P<0,VP;\LUAE[4#N@A[e\(JD[e
Xc9[O/H,?Ua<J,,KIW3@BS4dJXVRA3DQ\_#M+LE@H)RQ^(gLVZTf/0U]]T#\#^@#
WIDYgV_XS25e9OcWJ&WfNI^AC>g-QR8.0IgZ@@Z.a?9O_@-J9;W.9Id?>XNe.=^O
GQ;\]OdHAE&L1HdZN+4(>dc9V+MZO)Q42DG=2VHYK@YY9J7c9Jb>TUQRE5)IdIV.
KePV^55?b2SQVJPN^[(Y3ZG?2,02Gd#(/]O<40HZ)c@-<AJ7&:SD@Q>0C7BJ8O:>
5TZL?&(78IXeBRO#d5BB\R86]9][I&IZ)E8^_ad1TLX-+#^_:.CdgUMP_\PDDe6)
=E3W6>JL#E--g=R=e520-AID>cFLe@<Q5TUE_=9cKZJ5b+LDZ44C0KJ5=T?KJ1Cg
<6,Pe?:)OV)?2a&4M058E1>_D7[#,@CX8f^:(AU8Eb;C1MJ6bc;F52W[KB,:^Y<H
185)KH,8PA^.<9,M\f2WV3R/W_^?>(U/H^VJ)5H.5)@P>UJ5(D>TebEEG820EX<e
QZ:YeB8^K7c1M;-2MD;AY\_IS/;L&;R^#:A1b(I^JK>Q+dHc9eKe2bXg4/Q])>50
85H+MK)?DK+)_)3HH]JJSJ4)2O.ZLJ2F9O&+D^Xd\>FJ+PQ#[f5F+<^6OFS&C[Y+
D.^<=1GW[d?&KJ7gf<ZAJMY1^US<UU-M1CK1-E=e(_[]O#c8.(VZ0A\C+E=4WXAJ
1>:NN8a&DQWAd6d(.IK)XVCSE)<EU&[eYf<:24gf\LZ^Lgc)2G,E&bM)=:C(UJ5M
C^1d:>[RaNGg_GJI=Tc6dgPG@X4[LI,5EM>]5cB4<:UecG&71VNMa0PVd;g#]0Fa
5_a([#-[XUbX(>2a.]a^WXDgGEe#Jec@g,b0X[RNOH[#f=INL(;M23^ZB,@<K=BA
dWAI75W6b,-RdMZ>1.;YZ;4Ggc.a4XY?X?BBMf;<ME6:a;8Uc,O_?00Z:6C:dA]O
FS]-;EYW(aee]_g^/XE\]dd1;40NV][HQD6SQ[4NUaJZAJ=CeN)4RFQ4XTe,UP6b
1U]XQMQ;54^\Y3#=R2+eUUeS;6;/E8O4>/d#FLaeQE/C7W^VC5A/3X5-:Q0<N^HS
,SQ,,=X#7[ZM25Aa9M/S_MU/V-[?V0dScV+:N<=YIg5WX@_BCdVKXWLTD,)L\bSK
R;L^g2KGfCEV(e_?gPPeYIE=A1?;8H,+<4cGJfgDNPB97F3bC5L;df>.M&OG2WB+
&eQa-0+9YI-6_Mee8_(Z@TaS]WP)aEG?ePZ^_GO6c/@V\UP4\6CZ.Ng1@gd&Q<_Z
Hf_Pe6NPZWAZ6.?Y95E9-BePOQ8SEZ<=T_&g,RfG1[#/1<g/Ygb4Q<U0)WT3,G;Q
dX=cL;3]2cBN;Icc8]D-GY>0#\GI=5++(V]M;^-;CRb?+EW/Wa9Eg8E5+3f1@@-,
Q/\Y(-[1?a3#=BLgSRV#5bX4<A)AJc+@S/FA1V\//,AA/L9eT@R\?CV9XULN94FU
3^P<c;PWO:\6+QU1UQ_DWJ@-G:H_eL7b94[X_CI9@]LSC@bP45@2^H^40N?CQX^7
@BX+Je^<QP7FKFbL#,\5=T;WQ+8OaSVV-4aQc4D(f9RA(g]D_4+MADB^B8S4f<E[
-NCg)#GbYC+H46(8D-GKTV01;^2De+&fZ?X^8[_+INOLVNYMOG@g;dN=[BR,)Z9S
gf@,Z.5)7(Q&;(O-;F;.OX40#J>:S2ZNLDZ<GC&^9(^][,d-;P^gfKc1I31@3fWb
N):f,82ENSNX?)J#dL6ZYV9U6f]^U<O-L)+,,7A59^MA[@#W4a90LM>G<?C(02R#
g,2OZ(?EF2K-P3>O4@&FEH[]Y:,d1>7<CLI(0BHRd-\EYDHf,a(^Q@O>=aV1?[B@
S,]OM3b.BI0^2UeZ:,^[FZ30c4UX_C#V[PTOW8c9^].6fPP.F19.RVQO&DAW^SD-
-EVFISR6PRRZg^cA/]6XZ4bBS/d@[R]Q>+RMN#P0W5T<(OI4<9dX)gB(c1=5),\Q
=aOHUI/KQG05/BC>80<:)-T1@e0DL.SQ>,OD^A__(NN(L9HT1_@+7F\<bFH3\E=_
gN(bJ,R\-HQ4T]G4[2@[b(;]S4gY;6M\X#3^=4Mb)Y=KMVO=M6-Y0U-KR_K/=37,
5YKS)NR4K=BS=P;dI,ePQVW>/6[Vc;0C2>?^,Y_:NMQXg=aga17QX15(=H=Y881>
WF+Xd,X-Oc9&N\H^JYLV;P\Q4ggLMb.W.4<#R)@Pc+EF.(E^39\B6U2cW>ZLO5YO
VP6U(9]RO82;f+?Yd?9)f7N.(W\00bg#8ZC0E32:RSJ:,?a=Z#(S.CaMFG0X;O\f
VbU3^78cC+#Yec5C<cEgF:&D/^&01CZKLQ@:)B_=If=2^U)_LDdZVeU)0,)GC]EC
HeP3C0/4F&(Y3d>V^:70Q74N_N8-3@^:?[LCf1ZVT^_,+X_+U>F#E,(H(fL8W?Q?
e\6VT#)gBMY#R+>DaMD1Qb6,@5ANdR9]OgCQ&+>UT897WaNWIPY(49KF^DQ8I[0L
V#=7]D9L[RH.#6fX-S(1?==6^M=EP;/T=VBS.RGKHYA>QTF5L5OgA-<)[;8L:ZeF
23T=J.ZPT>/f6a4G0_F>[5QEffMY,R9RfABbY=157Z:-::J1RTXSVW?E5P,XW/95
b;H4;d-XET#HEXVK;_IG:@g8-GBCQ]4XA/F-D[bg_\NIc^,8&YJP3AV.(P,Y604&
&VJRQGV>E@Rb:;>[]8SE<N)F-JMab&EX]FfXd?\V991-MX2OQA)UW\L7>W7VTR#1
Z\=SH0@L01#ZI=fT@^f>BU?>L9S\JQ0a-ONJZ@T_OQK>3:GaWC0,(5_[RZcSFb>[
fQ;S&Q;(>=gBV81(g,,d>1;;/RcP>G6KfB9fPeC^8/]4bS.[7Z(WPB0YMG3(XgcT
REEU7X+E@WOGDW\T(F,P39)g[BG(S>)JMP=R#<;&cgLUbX4\>:cfAS<DS4b[74Ve
5NM(NNSg=R+O4NdA#QN?Rag?((cY)8L<abeEN/BY[JZ5T#WX1f=/.^\IB<+cL1e7
VHa+Y(aI\.1N.B,<J9835TV11O)67:UK1TA[48f/#e&KI;7RYWQ9YFL]&CM.>#3/
NS0:RO1QHdK<.g.W)d]VM+Q2b1&_)&b3U.R],>XQa?=a3a2b_\-;]0I2[WK^9D(3
dBFF(_?07G6fQU<23R)?;FbF?>@P-I[a;DAOKeLBL4-C\]KZ+cC]]D_:CT7V.AT=
c6EPZJHKP-:I9EA,9:\Y16WK,?J8:R\A-OF>3VYR8:<)BXd58/YM&?@#V&OL&<UY
D2ULVG-XM8J+:9U=)8bHI(I(PB93e6JMT):R5<3)YeY:c@;6[cJUCP;1.485G+IR
T3(^Ia1NW;-E/aXeL2AdDKS5I>Q#70@,9.+PdI_/=XMRFCOZI,SUI:EO-R)8gCM&
M_9#f,TP8gDODYTM0.Ng[0S[\E=ScA+A8a-8Y_D3NNJ62\:/>8UW+87c((2>cA;:
Gbag&@^QHg08ef)DVDQ8DRE2;[AB)e/44e-]&aRb2cUeZ[#cLWb/VVY0JJP+^ALK
)fCcQ11++19;)]Y[?g[Z#&C?K<IZD&-,MY#0D[,H]NaYE)2<VT@\:XW1dbO+M4XK
ZJ=FD[6W/6gPBf58_6[N\7-+J>c=I>6]b8UG7c(1O)d).YC4a36/CK-\(JWW:;.g
2GFA4R^CF,(<[>\YIe/4-fYH:UaJWLafGa[E10PE\OYg\1I9/G3Ib>GMd?^.=INU
Z3FJg3Q(5[,HCFPK77=S(8E].?FeFU,ff60H6PbfY;>gJAfga+3HdUcIE9AH59d@
G9//9K53Gg1Sf=Y]&QJY-W,@R;BB/2S5-XUb2,7,dMA@)YG9[5BJf?<;4L>VDeQV
Z\d/c;JAeFQ_#&^;bKP9W#.JIH4RX_T\P/01V37+&#9Ad-A>a3V#d&BGF]91X>/H
H7=\\2TUAR]HC)(M\4e<OeScHHW-4^:#9&S7_X_JA@;<gaY5YA);g]^8B\Qc52Xd
:XKJ(gVg2<43540A^@UcN6T/98@#)?I[,_BG1ED1#X^WgVcB)AMM8/\,d2WI^7<A
b0DYM;Mgb04PJ]BCGe?^R;J1-I5Yd^YfB(N36&gBZ,U7Z8LPIe\UL)5=SR]eHO[8
M)CM+71J_Y/T3-/XY@1NQY&,+TEF(EX95&0=;\;8b4=\LX1;QTAX4KO+GI7fQ5f&
a>@g0]N#E(8<0NUMGbOg7AY\)fONCU#QD_BP67[dA5/d_,92]gFbBFf5,0#Qe\I1
K0a[RV7,C_6+<=72EE?QTgAA.2^GW]eCPN&2#0SgADB=R\B;7db@&EG(PfI]<H>;
5+/g]S[F3M2&W1a_<B9ZZ-3;LJU504&;fF<e>gDF[?<VV.4K4/La;W2B\T;D9=Y9
6^V3ced,/>(I.4WNJL9I@NM?3N11,[.]gf;A+ff,?+LWT-XOALKbI3eeK9:dP_(:
NVF:LWEc9&@LX:G=Ac1b1H#11,)Y_Z2Ie\-8<^PCMLD\/Tf8J/&W[g0V<OGZN81/
9<fAUVZ?caXY?V?cJTbJO(>bTE(MJ4U4[Z?-?\4;X(;M,SeH^d]P&5M)>-G]b63.
IY[6^6XIab74Ud/0KMA1eQ;eD/HEF,7ga#+?JD0FfQD(XW-(ILgFC+bL7JdU/K)D
^(WB4>cHND4LDOB-@bP2^Q.c]@?Wa_(?J7EadEG^6V.0A&+7dP[4\M[bSJ[gY^,c
Z,J+##8K_[?B&-a#_HAa>7a3GUaNNGd,>:_H@KH1_M1gX-7a6\a,I#^L?.@[@G;d
BfOZ^]gTed6A_ST<MVPB/4MJ-]JfRI(g(Ja2KUGKX;.-<.F55/W4/@&Tc>0[6D?B
4OeeaO0gd6ISVdW]53.#G5,IE=#NHGN^d&]Ze-TWGE)L,8FgIE2H]H)dR_da9FV4
D/7XQgK;F2)8M.fLFZbO]5P&7(GQTLg<9,7836#ZbL2dW3O4V]L@2Ea5S<)+g?9f
U)f<42METLOEfX0&;OPfQMS>@9P)@?#,6Vd]84KP3>aC]9==1A@3bPVM,MI6)E<E
UO;EX@)M18@B//5Y-If-?B2dLd1WUV_6)B:W]+PZ8bIX-YAVVP[Dc<:H&\^cL44f
5)XedbR7E^K_VN8/b6+g:(W<+CdI66a:VX.&FRM9=2:>>R#\T1;IU9IW/VU_J5Y0
3d&#AXe1Xf[ec8SPC7aW=9FK>.&RH)Ra/ILXGZ:[Rc[^G+>1E?GTL^(6+7f&:;5[
)D\21F3bJ7/ZV<L1^L+dfe__?c>1>P6-a-YLDD;^cR-b.P_B6@4#P\MRG1L?\ggO
6G6a)()^^g&>H\X#(VR)0)ScCX[KW+,UK[)>DUXSg,QcXG]5Q/FO[dUE[f7;c^VA
DVN3cfHHFf2N2[aEd,14WP]?)6bb4&G2+g)9UeK>(DT/+NXA7,)L?0S&23)2H=JC
fUIL:-T5IUCfEY8>cC-)4?EOKU^2KSdc@T[.Sf<S@8=f4>)79<@[H0d(<[A1?+49
7)0O>T0/?BN&]R4&a3Q\bJ[4M]4f)bUddG@[?YbC0E=O8fC2OX3GH6./+)QK.^#[
c49[T]PZgMg5P<d_A@;?J4NJJS0:0F<,&GZ>;:/QdYg.=IOW,Iaf_K^TV^O1.d;C
S9XSe#7RNJ5f,2P4&&14)]L1eg4fEKb2Ue_eL(fOQH=R.SONPAdY3QQP&N3a/OVW
P0Ta+<9-N+0^fS>8(?1<O,[T)6/7E8.OY6BAYI\.4gY2;fYEH?,V@YaABKG8J[]b
&ARde><NSWfIGD_UGcb,PVf?NaROd;/9\F4JHLS_e+Z#1154#RXY6FY[JP@2,M41
gAL[\UM)Jf/U^I]E:AN3^1Nf3U\ZM+[LKN;@+Fa_B#GUYB.)+BWd2Y>#LH^2<K;.
UV1f_eRYg5#2+MReFJW-9EQI@&-R79e/))DVJdL]LAKQ(:eS>)3Z(]QeY-e3IVOM
;@-eJbKK][Y8R0eUb34K3;W+PX,FN-L[@#7=c&V2bY#0);Y)f?Yc3L7Ic5Q0HHM1
+Q-.@;N>B.:T7CNO7e)ZW=\F,Of1Y7<MZg\QM\b;34S3X?FH+,9a9LZea==Eg,+N
-FQg@3@=R_]T[8_5BB4\6G8C\-^]7@QFAS6TUA?Kg/R?ST:L>M6/U[Ag2OB/0M<1
M9<,Y@.?>He1a_-@ACbG0NGPVFG+?AFM-=UC5M,]e/R/9GDOb89Yg+#Hf2\fgNJR
Y3cS=,WX2;UO.#O]gZT0QF2>Q8ecP:D:&7V50^Ib5#J/E;Ea55bW]K(XX4&0#FeR
EK&fF?e)^FI1GO_DUE-?C+]V?M9LgZL/eHM^I,]eK^S&IgMT8Q/Q99,+SOPAZG6N
<XIAHOD8(,F^Lf/CdQ^5:06ZD0>Ga>gOd=A#.:BDOaZ37NOZ0[gD]8M?&?6CD>)3
C9dD?J_U[Nd55Q)[+548dXMFZ]^3NC9YH.W;XRM<08aP#JJ#H6,,@+OJ0K]P,F64
fc\;GfI@,_3F+16J.+Cg_8a0,bT[4OFCA6H+)(YSP@&GGT6)>U.-(19E?cG0]<;1
U)2[+I;cQ<Q^_RcF9/LbGY/48Jd8P,6XSee,8(PF?ac_,WTfM=K_CLaL;2TJGIZf
&fW2Y^_?2&.PW7fFaCa86ac)N(J>5V@Ma:81YB@>^Uf[-DV&MF)WdWT^=1B;,FJ)
N=Q^6AWA.TUW+-?DeM,J1TdMaDIE-@10B92G=C6H/\YEL02d^bX2U;OA=dX?=/QR
AVCKA4,f0C8@d5>#OQ-3FAEW#MfD-\X=5Oa;YX9[JJOE?WKL]CWL@JBG5(90Xb#e
8=TPZc:D>c0(&\G4^W=\W3^=+^<GUdV7d.):^)5B4?XaSD@E<^QW[G;8dM#F#X<>
VbfENRVVA94^Va,C(OF5^Z:&OH8G9e(a+RQC;(1Q5bTcWLO3>bA\+5A6Q(WS.HRZ
:30J-SI1>_#QT,&F\P^BI5E6XTd)?M&_@]W#:-M<76+Pd=24DJ3M9=MY7&.68[TT
DN<4]HCb_&1PFe0NQ64TUE3#6//X1fa2Z\U;@K+TA.N^]05PH37LQGCX6H7A&5=G
)TaC3KW2P[KG16Q+5]IYb](fNM8Q.V4N,V,0Z3gU0]AcRBD_L6[?KO>3TJ.W9Uf1
aJJL-+aC;O-HUe\=RYJH:3<(_g[Y[f]:?eQU.<U7T::P0If(Z=Bdg)J^b)40=\#K
(&<3UJ?>N.5[CFHT846B@S1HMZ<Q5FL9I2RZM=d.FF@178R/DONGVgP::0aE/@NO
/QBLV,bGf7_0B-c\Q=9>O#0[aHX0#?2g:X#B-YLIG.(:fdf-P-.3We@J>#/&@<^[
G\Ic)<CR1Y=f1fb]Q@T:O?Z/Q++X\\g?(a@\]>a2AY3T&34aHDI#5M]#<d\M633A
5H]&8W9PO[0R^e&ESM57)GWTN-<D8Dcg\[bS1//5\BJFD]cfJ.)8=FV(N&9?@V,a
E=GOX9T^g81g=[;4X(7O7K,BLUTS-,e1(A/;V+JIAeeT[,T2GbBXR+d@bH9#-Ha@
(+c6,D9Q4_J[1JDMa<]fO_EEIXE8a]DXVRK]M^1TIA,9G_Y5P>?@FY<>(=0>c>05
fDXS@8FNEPS^AZV-)5CcV8_LUOU/156bAgd=g_[/[dVIb8SL6g9Sc<6J]VRCHG<0
)^1-:g0&Q/O1Z8NNW[E(L(/gcV=HM]ccMS9b4V>V._P;/#[]#IT&.\_KLCUB5ACU
&JacEU@LD:4AK=;@P8eWX:[,POW?:S2?+0GQ^ONXC)D<Bd8JS)@F&[J:UN3K-9</
-gP-23^O/.)55E,eNE4VI]BZb]1b[+M.fARM(=A1)+=2H&<-a(_3\>W:-T(/_8/M
D-CAUE^<S5^I+^M](2@G-H58.#,bc?XDfGDO[_?>;4b=T][<LBR-76??>PfFf/ZF
RY)SXB1AHBfJO_V3KBA^1V77Ad2G<ZN>Z_Ic:d)1=#.)#9C-4N\[-()CHZKM7g:6
SLG?@f,M^UN-4XUf3H6OK1OF1cf>g^OD/.L0QUA+:X2ROQ/F^ffJQLS&Acae?Wfg
d6/PV@5eY>?EdJ)@f\\&7b[E+R@3MMOEd9B&YZ]IN7:G6[04_6^BE,WBQ<E)OD5T
#[7OOeB[6Q^,d=D,G^]:.ZS<J66AQ/_^N3WN:HKgg=/.\PdI(RG>+K\)d(9E]MY2
X;g<AGYcbgHFS1FAUg_TPG)VaP_XRD,[KLb.X:g?TO)<fGOGKT#-4T8Y)JQW+F?3
D6(F^KLVTO]1]R(ORT,W],4Z^&OZSLDXg[OEZ?M+)&44ZJ=&DcZ)O6@;KYQ/2>F3
PT]=8Dd^R9.CgMLDgL-8^1O:62Ed^7)fC.b:JLY(UGIWNGSOZMU=,SZ_W.Q0)G0U
^BV)0c(?87<<0OIf&?VFX=P9=g^Ld<fe[G<:_Ped85f[6Ef>H=)\1^(RU#(A8Od]
(?R^&IERf9C#<5V,bU6XDRf3_EeU#?;1;^/QH>H2+Y_38AA^]Og@+eYLgR3L@O8S
N@E=TP<cTZ5NPab23aA_&XF(_@9S6L[0&dOHL\E@LJ>X@6Z5L7>cLffQNF-(0eL-
e9TURHcD[X[bR=@QN_E),5\81cD;(-ZVFcD\Tc,5&MJCbX-9ACB<GYWE;8(&g_L3
eI.N&HdOW,GLYbY5[9WM9HI&DA@LW9e8W-2I[N7^8DM.SFB_N]?G^<]\\E?[14K8
D=X_ON(+Sa#AZR9cZ1.#K0^@bZf#e.W2fd[=&/fHW=_DVYK0)8::bK<[^-g\JFN4
,+@QQJ^MART_4_gQ5)H+ERbX]C=D_P\O8VXY2Y&;d[@ef?W:)Mc71U;Z6?4VWXB\
RI;[\?,eg--ed(\85MG?R_EBFSDF/a_[0=)<JGOgO=8M#bgVK<??EU4)@e&IbS;3
A)U\7@:Rf/V3B&GJ?)?GN<<AAfQd8HLC/YUU.;a7Y:F@_T-b]@N(>_UVX&RJ0BEa
9Z@;3\&?S-B;-f.C\/^.#bTQ)@NUab7#^=Gc<g&.1QDQ53,B7>cB:<Be_28@eL45
KWa2Jg]Q+?;85IR#cbEFZ+((geE.R41K#&+8e:[-/KEFH_+WU\7<R,7PB:6b>B>:
G9@VC0,a]);F3,BYH3DX39U<Ca8IWgLc[1Y7+\)I.TUACV8,=Y>;I7MF1T2._?X.
_8]#)3VRPHQ2:JB[7B.)cH4R?F_?IU9TT>@d2;.7^RS2PT,I9E]2YC3^+EBYJ=[H
R,G]A.PN/I)E/U^Oc,c[:fb0EI0])K-:CXH289XWH=>3B0SK78J9F1a3_R21@^T^
-:0K]LQX78?1PPJ>R=Qa,;A:\]g=<DUd5FSK@OV&fLD.6OG/8g_IV3-L?YPFHfL(
;gA;eW4[d4J?d?a@DN0TG]+KD3GZBK99A8)]:HV_AgNN]C4;H8]S523a_0@c7V2?
3W\QMe^U76<c2FB4\Q[53[ODaR2C2(N=a0XIdCG6(PYXGG)G<g>ILOVaLUJ(.8&9
be4TNf]AT6^^\2g>f,-2Q/TJ0:->Sa?#P)810#7^&0I&aD](_CD<_NFf,\##4_=1
g^0(:U6EbR.T]KOO=S_:W-YEgJfcVARQRLME_;3=Y0E+[54d#gb,M-OQG<6&>(CL
_[=Z_3([8D^c9F(I2-9G&;1Y4WV4?\aGbDG47>(9NN6Z,Q-gK1P6D0#JS8B5g?PG
97(.8aE\FT^KHOe1Y5g>MW36V,WLWeV>ZF\6];.g;C/D8G1eI01PDD..La0@L9b8
O9A99^52TGWF0cF1(?7V;_URNW1A)4\HdbWK[A2d@^9]50E2UR?&eb)3JS_a,\QY
Z9T2LW#X^K0<N;NT/#B5W86CPI)+UD7TWR5IX@6#(,]CKO8)S&?7HEg.3H8GXDOT
[Ub,fBK)OKXT]7fdD@2.O#2gZbNId=Td5.3L-C^gRM1].Q0c(@M4W1b12XD^@a5:
&c=X42.]NDW6d=C))R?8N,e2),0.<VdK#O&G6fXZbW-a2N(Q5LE-7bJ=@].eK?d?
+aBc]GW/T>VMKcMM.VR8[2V8]_8=[)QefS7RXR4QE_)+/ZX>?B\YD=^e?TE>/gb-
#>(2RZ&DG0(/@AP3gX-aP/,OaL+_A^VPK@DSD.=<1(BRNSVLK8[PO?[NdO,6:X:d
P0]W5P)[@;C7D\^E-bKb3X>(fB/>+P(Z@XI38d]7eGP@UY0Gc>OFQ-)JWHV>eE(b
_bcZ^OR<^a6W[Y4)dA\?<P.E=.-2TX)1^(RQ_-a0O3+eTB-H3dDD^ed<7S@>8T_^
/Of,9JPZ9BPb^KBAK6BWNH;[=]1YQ1R83/TE,UW7KAI4d5<Xd;:G/KX)Wg6-,)N>
2AOJKIZ-(&]1BF]_+\BKdd04_4=/(^^MFb[.--0=7@AgO0@eaGMU_D1REILJID07
c.dSR)[60X-X4+6_Z_7Md1D-JY#FLD6?KS+IT->UW)Q(0A..G8RN?1G@QSE^YE4F
\EdbV65_gA[<+g?DGK^-cAbC\+4&>7?L/YZ7?JK037CB^3YbDg[]JZcQ+<EEaaSZ
RD(e3\U>MRRL);+Q74Ne&)E(.I0+Nbf-b_X[M]ZLXD#?S;;fgIK6L#dLa4f=6N:5
;Za6[Y/U7L(JMfQ[AUPH1(BH7R>4Q:W.&VQA>ea83=5+W>AE6>]DfUP:BEVOc+2[
CbCa;,0=@^(E#43Yf,&e1,ZC0/-1S(=CC-Sc=NRaeB/75R2@NT70XB:cW?VP9?)H
)_2/:=AN<KRcK-2HKIU.3G^28N8XG[_ID2:#_JdcV+81<P_Z@e/6_>F/-aRM:3^G
3]d_RDX1>Q9?L,F5WTN8<f+6[8A23bQZXNYCUcNTQ930U@)R#a2J;=./_d.N#31N
dH,^a:+K@^A9Q@CQVc<^2;L66M\VU.T;_7g]+3]\=]JA-ZB.0W.WgRK^;I&,E,C@
MIQ1NQ@\<-B)JOWCfEB71IHM07Z&HMHP@QW>+VL1OGU34XOUMLN.M?B12G)GD#T[
D=F(aZ>Q?+VaPXYO([/03;WDZV;(DPaa\>-gD_I&SE/61,g]EZPA^\?+F<9>R74g
T^^XVNGQT&71ad7L(b1:)M(3@+#++W66CU0Y/_5SdJM0bNJ=de\G&;95XdBCbJOg
6gM@]M=@8e7W8Ze<a#c94]?T9VLI/CFca=2;4TgCOAC^6+Ba2_NU=S-d[4?7<UHS
6;UY[#4WN\6[cS7Y4bO(0(9e_VeO_)/OP4.5QaK><HNVH1\HGA:E#a(74RU)6DAf
[?3>(2-\/D]NADc5@g6RLFE+6CJ>CP+8a/T;G600?U(M<T^EKcUEcfeID#a279BO
;LFO6c>-_F+OVZc<(fA+LH&G<:X?)K)DEG7MgJUA;P5C2J9L9#[0dAQA8IMY162U
_T58U5?R]BcJ^GG?UHg\H5YV&5.V[;8DZG/_SH[3fP7BMQQ>HaKIILEDdL0-c5;&
7@(LUA9_T:W>-8=gJ([2=U?e)C-3,#.Q:B,>JA8NB7Y]?Q7JgMeU@E5VcAd:WRNN
Qd>]/S^[QY2F6?>c68B/3,;:&N7/OVQ>UBAQ,+=a+Da-P3Uc_^^LC5WeYNg/.F0@
[d\[GU^ENb_4Nf>3-]&CXC2?S5CU05Id5Z8J1J>Gc2NYdC.EXfM>M0_NR/\7bF^\
gK>>KTN-CLB;JL)&3cQ>IX0N(K/T,:cEBS12B;2cKU.^T[M7.OLI]#6Y&IQITUMC
KG><>bT6B1\7N&/X+C1fWE0:#ZI]]Z6DQ^:FR&S=0\P@8+GM,9P&)<8214?RI0HD
[);6Q1HX><)/,FFM./5@__WZ])bOD1^O&E=7dIF(G(BQ83Ub5B2N4\[K.9O]AD/M
@d?HHPFM^VF/)$
`endprotected
