// `include "../00_TESTBED/pseudo_DRAM.sv"
`include "Usertype.sv"

`define PATNUM  5400
`define SEED 5487
`define CYCLE_TIME 5.6

program automatic PATTERN(input clk, INF.PATTERN inf);

`protected
;T(d[VTg?TcNd/WZ5)\[ARJGb&(LP-(=1SMF.e2GUZcD@UM;C&>I3)&g1#+[LRT>
;F(=(6V3;QV^Beg?4E&L]0>),INf@_+Q:()]a)820ZCK[dNHX0#TTD_,E4AXLTf+
ce?Na+?5PD)P0fJAQKXL9:KgN-V):ZW8AHVKV2YA_;Pf36IJ49S77Yb6TOL15,4]
2I5GDY7K_\D,MOf;\)(Z4/?7O/,W:@[^R=NZ;CQ[0)],&+C#gRH_dfGgBQX]B=IX
IEP2cMXTE^7b;VXfa--<4NLe3RB-8@@(N;7aCANW=Cb_T:7DDJO&d&3(/R6_86B9
T,^Z#1(_d;J9d2&6YfF:4<Y[7QOJ6LB\Kg:V-eY;2GY-\S:bJU0[/H3QT@XC/)<L
7aP+A#/3C<#5\R,Ab2D5]f<RR>d6,eb)1R2gZF/<R0E6#-(7)6>G<1ZVf^T]F#:1
g03;F&Z,gF-@Z@<McZ8S.B@Za\eZ4RA]f2De^9CF(5.YS,9P2(ZS?IfR68H0UM/V
)e<<19L&Za=]XH5VUA59Z==EU7F_e.\6b>:W\NE77/)c=f-M58aO4e-YXcS<:-\=
X[0XB5bMcg<5C=EgLbJ^O(-g)LG&?.;J7GDKb48A&C?Db8J:]-.-Oa;B96))A7D7
>RYZ(gFb\aa>Z;,<c.dPACSZ,b]6]K3+I(.RgH(E:(?NCEBG_Q^8K0WY]4+BTT#]
2#.Se<=YMDW2:\;b&0Q6&88)(C\T;TRUKe]Of/FI]7T39LGD^C1L3&?@g^?JBX]I
fUH,6>DQ1[Hb@XYEA54-&[=779Y9W_g+LAZ\+BX6d:IE)2M=C/_=Z0N003d<&&W8
M[F6V@@-=OFeXRdCZ_X>L6:N:BgYY)LKXa],aLFe,LEW(3M)[b,61L4.6CHH^1Rb
a)A=8aeJWI#0+:fcdfRTS.7@JBUV>41S-DCA8M+?dNfP65ERbT2/W:X,=,+=F:LG
64)bN@>AEDf:B@aP9K<-NED5:Q9ZN=9A^O7XT?Z--6^B]Y1_,9FDfEP/Y4Y+PU22
BIcFJ;-8K#g7)W>MEBA)W[AI[Z1.b_\f0=CN+&E_L3>55QBE^D>=eFHIRF^YQUQ1
,E=:b]DDfE7[LPLUg.WXTba&3,T&@F<;8F:Za[Yb2^&&EM]/Qa6C/cPW7F=KUR@X
G2:EL+HVbHa(6MEd:[.bR&Y8J7T^BJ+<E3ca9<?f5M@Bf^0N43)_aT[96W9X?/bD
M)F-@e4Ff/079Ab3[62GIH7^>-,7]=1/6P/NbFg](2.3T2Wd6I,^eX:(c+cVBe-Z
;)gKFZ6IX1b?2+<)#PLJ313UQM/Y].BN2>dg<1\5^@<2UF=CGA#5XaF4C:7&46^;
B\W54#G;U4d1f.JDgbES))YYW4d2a@@<>W[.0g2PbDdZAebQ<8b>X>GEfXPK-I(8
WS5/?OC=L&B6G^W6\09+a_cT#\?_PAK1GJH&.L=QV.AHLLe_5Z6+CIYOd-7R&]aW
,AST_EB:?[#WF@H(Y@?c8bW.9VBYXCX;REBWWKPef<&/_0>GaL#4-5LKV>FWg)&7
>HOR,G1WA@AT-U&5+REe^#CeQW_GP\KXR/T5T4>ILX<W;2;=JZ_B&(3.]@<N98Z4
^<_X)fK&E.A1;^ASM)T8)A&6U9(R7bb.6I<#,+95SMcc)+BT6E<Y\QZUA;S>3^P]
4.-):8M3,@TCZ?Zad/,X#;D)TIL1)IOHU^OWc=?gFdDJMJJdY.[#)>UHbf8G3HT:
SMcT7aNcfaJc[:>[4:GE/?Lb112I5YGc_RRHF70+_?8>a)=&-^BBMMgA[=;HLWMW
3)B6U9);]0)CPSE?T&A4af>a;3B4Nd)CXP>We(U82feZ++V,7W&F<E]dMB5D\Kf2
X]75JR3dQ][H-\\+0PXO_0]N/Ig:-H6f&.8L^.Oa)WQFAGLCJ@5=U<4d[0U:MI6\
3ef5gI8U_V@=02J:JNZ?Sgcc9RB&GGVKE8UAV4G;MEWKHO^f:;V8A[,;J)ARGUFZ
d-S]9X2371\&@,D?g,N+gX3FHWAI6fGe_;f=EB1SL0Nef?1>NZVaGLXH,Xde&H^e
HK^.Y@.3<7WP0/<gKI4\VA>/=O\/6^#Ae61@GfHM,Je=QL,2UT+:_03LV)gDX.]5
=YaW3U_cC--e]\GZ@#E\EAH8S7F@d>NFTM)01f<\7A/0R]0P:Cf^_aS-&bY51d,+
.P0,E.f?9;;AI/GHg+^#20EI@gK0B][R-NY1K)XdB6c;cME[,AfAT(QTf3?PA7UN
QVH7(-B1>?@.+>O+9J;S?ff;B>MHZPNgF)L:AU<6Z@>332&P>FdVLb7c@VFM3f=P
8M+8G4XQ?;dXSe^;SEI#3_Ea?FR/BC4L#\@,&)DR;a[^G[BH:SebQPe_11HF9:UQ
CZCMf\5:KUZg?Ncb-6(S0-IB<9N_R=CO(7V#WWfS[,Z_83NOUa(?Q?CG_g#^WB1W
W;OQPL#[,<0G#f2B/K[WSRNc0#F2UYQKE-S96DVUUS.UF,<4\63a-1_-SD\Q,>OS
AfUO+b]B[^3&([d(^-OB@NWLf<L<F&\=2V&4(DUC5d=&:/e\.9FX3+,E)R^VE._^
664\W\H[SUc?IVbPc5YF]-:;7I2S>N?;U]a;#)a[>5LW6QT8=6R+16)]R6-K^GGC
gd]6X.V9bIG1a=]H6F.G5O4>HSab&8A)BWcE<8ceb,+/X0OI9,FYgAE?8+0Tf7@D
Q8-B.+A0,8g&=MMZK46Fd4MXCIF,&RBc__1-A]:I[PK=MOb,/?Q,T.4-FRe(S&]V
\=2M#5\U&D&[)+#^6_IHdeRJ6A0U+A5be5a3gZe)PHU21)Y#52TH-7PaQRDD,V25
c7JE;cgbB\6S?g51##/=2?-72H@-##MV[O1dUC4533,X/[<BX:a.DcFc8V#+M2Jc
2H?O(^3=II&.-EDM<1.8?8GA2Ace6KL]DRO0=^TJWIRD\7aIA.Rd+\O1[X+TMK6T
30GFILUL8+;(8+YQga/DX,]YV/EF7b+9PfT.AIC5W&?S+\ZGT9&+f3egYPJ;U@QE
a7]YfGR3H1bUF[MB2[WF.H9B;[#U>;VQ?5&PV-8TKC^P:Je)RAV)ZJLfF8KXgI?L
g?,(ZggVV#P,-PE&/8W&/PAF3SB)>=&>NLSOf:(Y1.&#0F,gBUN5cXEge:--a.P4
#G>gJfP#?5=,UNN7MQgQId\7YbbH3P8#Td46N,GadbL5HG43>MLGU6?PfG6M&U4=
GcM7WAFTQ<3eV1;BS@ceUL.&CAID2GME97HJ>IOT&TSKT1;DP.WG5YGe/[ZZ4<<5
;:;NXgQSW+#U-X(O^5@Y4G+Ma@5^.:HJ[1EA;R/_d825Z,>4ZY,/Z3X&\,?7_M_a
&&e4[,T;15E,FQe96FL.5JeVT\-ZV_EgG,E,@L.,EJ.32C.N\=_LQ@)>NH2S_&bO
)a>?(0cNZg6VCaWQD>f?^]ZYGf+7X7Q&]6T^^M2;Gc;b0b2YKFNOMC(X@QN_g/NY
E/Ab,88XRGNc6ZS#J,S-_]_D9a:2A7#6P)NJ5I)=M-3^.6Z;TCP5-EZ)JE;H&b-K
U9RXd8A;aN0?0eM1)Id(ZQS<K)J^QDHTLa6_B,9RCID:6BFWc[cLEMVf@:\49RH3
#Taa6+D;<@<>-a]U?2:-:.<8)+PBe&AK^?<_)RZW25?X:97J=P0KZ-XJ.J>^4:=M
==@Yg44H>.-)bN/RAF?La=IKa13#Y^0+[YQ&4XWL3BI(+QKfJNL/S&,J+3aCA8[Q
9dfQYV)#VdU5L7)?Z;Nccc416gGI(NB4_T^:Sc15[\_fMb=Z[1WQRQOF=Y;4<\>c
((dg:D#(A@Z=JK501=3XTT5E0WBLQH^=B:+[]D&2IEAfEBUF=4-eIKQ:09>RM]U]
1aM._IAL0>>=>R:;(=KCID9/Q?]ENI[fS0C;P]7NC>/\KJ#O.f.GeeD(?X#1BZ^(
Z.RAZKKV_B4,,fW/^EOKAea3.ea@aIDI#fc/PZaR7WfK9)bdeK<YNdC2+I0C@A/G
[dV>#U(;L7]?,gMbC?f<T-XGA,dP980+\[^8R-40MDR=BK,e]bf0<@3-QK1E(#=1
gKH@?X=eg@0A.[N(^-T0>G?2S_880XT#HLNVU,T\OPc6#\7-D316NA0)DT_-Ig6U
d-Nf>PSF8K0:KK7\03EI0G5DW]27#27U0aS[G[Yd9)7F=Z[AC9BZ8X[F33&/8\IL
,D6&5-O((]WILaE.dX:J?1XW7P@/957XG+#G,DP3ZTgF,[ELJ++<;^49=^-F&K^3
>2gZC=,-YQR]Wc)TJO\NIgN:a83]2H]Q5.]Y=&:F]-cEf=cIdP^=@([cQD74e10O
f6NFa?=&-6UMcG8E:V2HIUC+ZP0(\=4c73,@@D3(UPMM/BSUUW?Ha>d9T;)22^<P
Ee<BE3\b//<=T?5F3[R)Ob6M[L9T,bfJ0g#]EOd+_G68(4@L?b&#;d8+1LCLOSHc
[R<]6:(#\^:cI>;DPN@OFdSBPQ_CKMV)OP5\.;Q+b8fg,EW95G:2gfaZ6Ka,AC0Y
>R:#YaP2Q;.,ff^bJ^S^,C3,0OV@T<0C-L0IM2@DXHW&-FVYE>I(Y9V1d?,W5C?E
:QQS_.(07GAO6Y3WBC4d)c/7\U[e(MJ6ON@Z&QO\6Y;Ff;,PWN;CECL945F126:Q
##X0HbPNPZfRABFeG0<d1f,XU&b9g_.6(>#Z;3OEHF?PHO7,Tc8-TBVETQ:[3.LI
9HI/e1H8.)[/PKBca,AED>;5@e^C55EgM?UKDPL_gaRIgT:<^F57W>3I?VM<a4QH
VYb5bd7EA[>M:2@P_d>C4?gZLdNMTa=8+:X=>\?P0PN4@HG)&2XP?LQ.EB0/JQ&Z
7Bg,-@8e</?--U#=5d?TZ736J5-]?Dg)9#]SNN#CA:GL<-91>>NAHR0_(9WPCUWQ
:),->KPg1G(2KCTI0^WL]d(]b;M8:4L594FY\fYa>B#N_8Nd(\7-0S+_9#8H2@g3
SQ#JbR_<YF12bE0-g+]8XVA+&F7YTZA\72/eQ&19<?._3N,7DGR4V?B+<<\5..4M
7Wc.]M_X]\bc;-M2a_Z]O.QD37H/)b)Kg^g<M-\gZ,Nc>\34A+R.f570AB9S370f
,PAdF-9BZfXL16^KCXaLRWb<ATAR8O0)D6IQP+V,WR=Q)ILRDZTf^]?,WQ6O[7+A
:e8D=dOTRO^M]\d=.T(D6^CS6Ff8T,b==c5#-CVVCCa3fTBM#b/1dIH5/<@2<A48
Ed@_OQbcPD<O6dO&R5,eX@\gN[U(3+D^J0;QI7&g#:>E]B2bLY-#AU3319_bZJCA
VL]#@>ON_,dL,b\V7O[/gEbFGdbBbdLcc9H^0d13[2f0QQc&9b?fDAI1<aY#D89&
VCNG=\faE9WO;.:Sa9.CNa4:OWA,C=EFNQe_<:[V^SMODf>7=C0.O#2f8SENTgVb
-I;G9+H(.+.8UKUP.[SY2^P#[Q\.X+<X#_7d6=-<GA:TT&4CQR6S45f9?PTbA2Y7
X]EH/X0=CXLQ.25#WN)2-Q,_@<ad\[D;-#a701R4S^72/J_MF&Y(&A29N,[-3OCD
N7.=;\2C6+_92AWJgJg4g>71@WdM0TSGJE&8;CE4VbYe@S,_9@a,A@Ja]<-D]5_6
I0X;4/#@NHWW309d(.E]\JSA@KBgY1(_IEA[U4g3d/e<\HK^Z9WQVH\RRCbf+dCW
?Dd:=)4RAJA.[M.g;XZ^Y1.PIb>/+BZ#d+I:[A.E<QfZ?QNfH^,Ke.NUHMD-Id2)
M)\_FR2YQC4:8UH@T[96]&5^-&-Ad;G=;K4UFK<[Q4agKMWB3,MY)fSQ?6c:XdHI
KBJ5DLET+7=b<:d4QK##U?E^BCNd0@KgNV28K6+^&BSHbSYaKYC/d9X;N/3I#PMK
e))H?G488?.dYCXR624)PXd,4=,#e0LYX5/LH8Q@Y1VSK4d?X+.J2WXd\4C.ag=<
QOKL+4+&P#LIN4&=G(Qc#P-.F0V]=FW/K];)2FKF>IEV1@adO#3#,I:RBE]F7+>K
V,ZY2SF>IRMaKZWTTY@T.@]S;][MRR\e29I2d<fdL[JHC3G>SQ<@O)?f88HE(9JN
NH<:0^8YU(6SZ2EPIW7(Y]1e7UcDN=8DYK0+eD>TZGB#5=MLWOIeX-5KH6J,d=U+
6UXQX[A2I)1Ue-P4b+YcWPYVG&/VL^GLKF0@)1^&=Xe]8gNV<36bP.@a^#baE>^D
27X28)Va(7WRFG)A\[[\3.@K2.G5/.Df9@gBM\gZW71IHVRYU^(NFYR/17X5e9Y9
:E[[cB+=R:)OT206UO,,RA.Z(;)R&K_cJV<[cZN[EQ(cdCVM]a\K/aC)ZB?g5.c-
,?:SaABERdf,X7=)<0bP=FELaU7[@7P[XB6_^/RAB-NLWQ(55;&4Xggd5dK6GXI>
Z?b^.+D293cQJ\P/5O,0Ia=acES,S[>#;VU4GHYXJX6@EZ9JG&WE?FaT<OcN1\E_
_T98Z4dD.0?;=D@RC]T4(3>7Q>35MP[4ITNU1H0PM-PWH4=B7VaSZ.SL(b4G,[@J
?Y873ZcKB.,&=7SeDa9JF86=e[>IH;8C\5TH>S/3<#QNUDKCX#H0AVV^&]0P-9:,
)\a/69,=E6/<a,eT:;eL^;Y8fA5eV4]Y4S6S16aH:,.E8,2-&VA1K:8d\0:8-HcO
KWWM2QfIfUKEV/_A,S395)c+YPOL:H_OPN/,)XH5f)\.[6B0;0IfI6fNA]BXf8HL
\.\=ea\NP5IEC,@)J/F8T\>.+@@REZ^OB1MAbW??[1L)G\,GW3FFN=]MU)7_/d84
O(1-7Y<5UHe?bZ6Mb:-XTTQW_C^MKcYd5)gSbfT4(SYN?+L3MOIQIJ.NV>1Y,;\g
gb?-@/L+1EZB3A=0&T?4I\(d>HGL.WRQ-LF:>.G8S6:K<cR>)E[M=GS?F-3C]>gM
fS=UC<eMO0b,JPBf7X2G8K=FgbHHM^/YX]7[aQ.gRL?P5ISV\-ZNA=Y[f[ENPE_^
II#Y]bIBPO-KH8XOO&#BPS]R49e:c@d17dXdb+Xc:FFB=.)PK/:8H]_49)c9c,N>
(MfN0L<0>N)65)@3abI()_#M,A0_3-VS-c:GeWJRI-#+<5<QcYaJa&XG;a9g3H??
JTKV]MU<LM64-QEc-e9GE=eIF9C,O2NX&Md,@02#AT+M\#EbS)?a[HE9(@H<5F?3
-(4\AaVWMS+)8ILfX9E/+.F(S>(]:;0+.3:a&b,2TgO:gQ:\1)H[72G;&ONMY)]L
(PD)[e_-IN2,[;K&;^2bLfcR@WPc3-YD.fZVWbL3MR0YO^>)&.SM5;<F,_T@4LcJ
.f(<cBD.H.GY@VL<E;EX[AI3TgX&C5fG<L>YT0>FENR:CEV7R&--Ld5aV=,J+@@7
5VYe<&Y_cbVB1FbY@A9dH;b4U7#_d=GN9@gMF--ZI-89C_^S-/6MPU;I;=:,<>>?
A</T9N8.aK6XXPLU\Kc,:CYKE:4dd(Q[-^#B7K^2<:YYW&)eAQ)Oe]If;@WG?-c2
X\Y,GOBAF1VeO85gf;R#LL?eHSgC6F^:58?9N+>=XX0N,6Sc,BCf_2(^;I=1g4P8
_SWW+K6/V)H->L/</bCOA.-M&LJOJ&WA+cQJ7:f>&YBARYAC_XD8\@@@bc2RDP+)
MCD.I)4Rbef,J,QHd+UM]+bAYX[M)VOUd+?M3K,J8g7P[dJV#HE9QZH#bf]YaGG[
>MSVOND>.e7]83(MIN^K=f6A+f;39(5OH&>_#1ZQ<9]0<F.7_H0@f^N#@[T4@(cG
;bd\Ng0ED:ZQ1f_L8,=@4ZMCWY>E<N1,eCa,7eEg#(7[/+@-fe\R/\YU?G/Q/g-R
N+Y<CWMM-OeH<BN-U+6E17=+M)FR^0QHP6U7-bd_3]M,)#AF&/O(0(b8f2L).Z,@
XK/B&6c@N.WH7]M1Xd8,^#6f94MI^W\C@RENW@0/CH/Z/eQ9UO0N;)\cS9c?OVUS
>2aA4-A_UE1-J](#/6+S#]+L2[[bda>KGPC5]X]M_,d/C<eZMX^GT\YZV,K6gDgX
RH]P9GgDcKFASAKSKI@:]-C^gJ7a+NMUR)b-fb+\g^HD26K4N/\e/YAfaW8fUW.R
]N]cgS<#GZOTg4JRH+GWe:-@YRZRU-g:713LgFC,0.23c,^V/4&\N1L;2I7>358]
B@G[8X[G&?]F;.-cMW2MFXDF_#C?C.GPT5A?B<[DD5;N#LTYY2U04GG35W256C5[
#VbHKTODMdf3a4a_+@0(M-&Cf40&O<^LBfCM>B2#gZgT;MfI7ZQN-e6<N:;WG]T@
;7S,Ae.(GWP-NG;+-#-1#X6/)]D1BN7M.WP:2TJ@97Z,Tb.5J/:eF<LW-.[S6@/O
)]+b0&1[>.^ILa8&bc@OE9D^WH0Sg[-LB;:g6&ZDYG,2Y@D@++d/.2G6MF-QC@G5
M&W73O.50V#.//g1N<_E#<YG7W\(.@:gf[-bTegG5GbR\Z27GA3VAF>?-JW8[F^A
=.I=\g8SR<_QMc52>bK@71])W)C/(cI5L(#ZVKT3&1VZZ+AMW#J]:+IQ]&A^.@:1
Z@]BGe<\\[f<=93ff;BJgY&197A1Y-+DUH(ZA&032RVR90BeL??XY/+=1[;dV5>6
.J<X=T3@bV,K>U;#>V].3((Fb_4cA0c[7)RIfac2+B2M.?8,65J6WE^/Q/K:[<P&
UQTU&>+W?8ZPP,D@)D>G3@6+MDFQ^Vb]8SRH^OHUc)NbA#>JS7A+0bSc.WR)7O5B
M@O)/DAW1eFB8IJ#&ADAVC&BG^@Q0[a<fX3\fd2>2#5Dg)b0ccQ-g\QX4L,V=(b3
3@RVe-#P+]UeWNK&GAD=KgLE^2]Me2:9Q4MZD35@5?/7[FA^E4g/CR+g#C2&2dTV
>J\TSOd=)I.T4>L3?9d044,g_QfCcC7;_^Z]N0,AdNDLFNeM@GW@0J;C][<c7\f9
]::(L60:O9RA??1Q<bgWdL((bWA)JgG^A;P(9Fd#3,S902M\DHAPPUT?d/)+SRET
3V8OE-,I4X2bHJe[9>4/=V.@A]a?EM.AX;MY,Zb4TU@WYPQd2/e\ab8)Sg&IC:,G
\f6[B<e>IQ47.7NJ5Od(Y=c-YbdKZgPQG)]21\IG1-6dAY6;R#OU:GTV7UEIMBF>
3b+(e;:9aY0(F_J)I2?ZT(O=MS:41LQ>g5_Ig.K7C99aXPLXe9I),HUIW[F[MNK6
be/\^Dd1KD/6VMI@6(,/X_21BSdBW?.0#0>35;Z<536S2QCaH#WLLF)gP-I1ASbf
)/IA5_,D3XJMF_IGWB#BMH[_IG5-O5aJ_#Ab?g9PHM3/M.7M.4ZR,50TP_OaQQb\
/e62CR?1B70c@#Wf]>eP,LHH;.87(dEQ5/((2K_d@)Uf?_/NM-QG(&^++I],)/QB
T=EgIGd&AWIgf<,Q5W<3>?/5-gR&6OZ(C_;CMI<?USfDb<Ab_B:,:a\<Z;7GHEU]
IB4JW)8?Kb:@KOVPJ2HTKcDOLRfNJ(gEN4C,9EfZ82=>6NNIDSTDf-C,-Sc2N4.A
IMYM4U_Q;TcELJK<=,]3>fDJB.FK3M\[9+W<)^U^dSdLOH@(4&25C\gNTWQ]H?&9
2gHDYbI6.KBM6g:A2Tf)La9:]7bA8fLYFDWG0SEG:#(]].SH,A+Xb(^9g.17WA@,
I5<,0Q:/9(TDHIVX1&OE7TRg(6b>SbL;[:dW;fCCV+VB=(SV=cS2Q^,gbT2a:KPP
-d2^_e(da@I;+SSFL<?VbK_L^g__b=VOf,LL+91O_A4N#TXHC)6+2;218TX@:,c<
K0_VMB0;ce9U;?VI)2X=g]8V<=I3,CP>YPYKX4A71===9P6;=,H[?WTC)W7B_]Q)
<8BB#TGP;L8NFSffCa.AbD3C),HE>/NEEYF;+@CFeSO-3Ae=8GNa4#:?F;(7N+1P
VKZ4g3^LHdXg\,XG99+4T0&e:bQK8K\0UO]0XN#2V0_ad25FQABf4GVNYAYH?.OB
/NaF>D)N_O\O()aX6UU&@-9:V#(NJM)58=/NaYSR9(Z6ZB[HXb52SD;)W+G249.,
-MASJ7^1@#5P#7/O8NO:Sg./2g,cSF(;,4M08;+ZN&(Eg3@4LIR:Y7-4JE/+<:M)
IQU1C@cT(LSEYX#I6GV7g1UR069gF,[1?e/@SA==CZ=[9dAO2K\Q)LT:ePNN)N3I
I7S13OH8/.(BIR)UZeBY\W:\a/4X@3J;=+7]1])fLaJHdK&#)Hd6B^MGGCCb..@7
)_E@G5WNU0EHb)UEZ(aH1M1gGI;8d6.Cc2COfJ5:6c2[2CC)S(_&De4B0H?L5J1g
<3c0.UG-Ne.[FGR5R[5fd:HSWC7>cYMMWF0^c&(<J+\5<c1e\Af;?OO3Y^X/WCRA
B+AZ&]Lg6&8^)DZ4U(KeC<>Eb)N;V&C=<=D6Z7J&Tadd@S/4<8\NE@/(:(7Qc2@P
#+[A>4UOT@GbPLg6daRfb@>X<CaT+/-1eJOHB@]>IBDAFXOGHMM,Ydf-_4.5-8E1
<\(9Q20W,#P/+_1K]=>2#aY4)N5;c]f/I+E,+XN/a/+P[E<OI_XTAQS9^+b^dOPG
7=G\/;Nc(QYZ&72:OF>&X5+TR)f/K#a5R5XTU]YQ+U9B/4O?Je=9<[O<XeP55Y=Z
4aWbP60L5#0.e,<79<24@GdT>65_FM_(&:b8/7ZVAXg@8FS85/=ET1Mb#..=YPL;
),N5W<>XJc>?XF<bd25QS-+bZ4\EW/b2BfYWA047DZQf\ZeL;N876eJH>1UE\?JZ
9]R<EfA7T@WQ+SRY^6Q<&03+NgB/_BIMfA=Z9H4-;7)#0WNWWS)[_)K/c6G/fJ57
g?QO])+V@=:P5H>LeP;.2b3RGDGYX_ZAL;;,\=O?305V+I>]PYNc@W95JZXBZgK)
5<f@FH)cB0Z)f?NV46f&c[[HGY4>P&#CdU-bMgX.3YY0I>VI>NRUb#QaMfK;C]K9
6e+7]7SH8^6?EFA)A)KbH&RGP9KP8T^M<0aW4f[RA@T65@FOT):)KJZ4LJ/3/U0J
d-5:Ld82,VKDeFT+-N=BGYAD0O<:Fd2N,Ke,XP[#275PK#a9C^BF]XUVRDTNL;JP
b#Na3/3(DAaS8HAgB9QLTFF+I02LFZ>3+@(XJPYHcQ.9FRS5-1AO,82XgEBa]6;=
ZL6I@<0f9:&^(Ue3d[R1g4=S#cE<JaX,Z.)=^8f0>Y3C9/4K+CR5UVL<]0BG&K6M
?,#QXbJa,6M=[&DdV6TY@b,#TJ34=9RfWQbOePXF8WJ]MBFF6U?_\J5;?(].PdAM
J]Aaf8(Q7Yca@,bB_3bg0bWI8D4+6=4affN1=_@3LCUZ18e>-Q3b-B+=^24IS<:R
@T_<?B?gLf]Fd8<\_EW>H48^Me(O4M.UM0ZO04c38BPD3UNVcGa1(/Y7fT1.I+/U
cI6@(ZbGCLLG0OZNAB-b&LGM5UBQ]f&H<0PZSK/.[Og:J7-ULT2OV/LDK<(5K8g4
1g.&\7[PT;0H7#cDC;2H#Y90PB:9#NATOGJ86a93W.@@L4RJL+E^gY5U,->A3,S>
U.c.L/8?U7\7I0CCDXFSO#c2\S#H9JaGAM-DGY@=F?HRRM<6H#Y6)?Q&P.HI[\8g
TW(OeCI-,W]f\T-=b,@)a@PLXbP/6^ccE;J:E/]CG;1RSNLdJ[Lf32)58YSS@AI#
]fO.M;AeE68UU)RQ?M#+9WL-;&_V,+eL9PBIM)b,RSBZN\VbA#P=<b7GB&P79PY]
25:^Z+8cF&b(=gRJ)P[1(E-5,?D@(K3G3\dL.,C3=WCEM8SeL3?^TIS,@-;dZbe5
R@gLd93WLP=J78J&g>J3g7P_aIN6=gd[8L.E/ab12FSbYRFW.7-LIbWRe]T7;,a;
@(C5=VeO9D/=2I@_JNVB0\eZ,/P_a,NHAX)/ZLF8)fRcgC<H1\.d?I]fGb_4EB4c
e-MI,\NTS<Ub2(3-9F#aL)2/5\Bd4M(:\.0;Y2K;fS4CY\bBVHEf#0_\)RL-&.cZ
7-#TP@+5+#c1B4Ng66AWX,f&P[FA?B2J#\GDIc^N;19ILg[3UNR<-6_:7=Z8VX=.
-fR&/?8^7H8PdC3VNJA:)-A>Rb/fWO44(599M2UfVdF+2N\4MT?g5V)cg]-RZB0&
d.NMUE0KG0;IS^\Hg[ASG3.45/VX\+BJ8c.E#TMY,Q-[0+N;cg[0_5c+ea\-_>KP
IVIC<d\WLLMI-J6GT]MNQ-O771ScA79Cd7=38b[SA=cXU+,==ENG8H,6GZ,8Xc?N
EDb<9(T)Q@AN2C4P\8=H(;,<HDKJU.fSWE(3Q=fFG;1LIagIG>dLg/8=3;J-S\KT
.R,cBTW&.0_[e])7Y#QK8YRgcg2Ff5^?Ic(A=D\BO/R/J>1Z(^)SXZLOY=edT<&,
]3X0RNg;d5&^DJ3Q8ID@Q9F84^3I,TcgO9b6deAB9)[MW,L3?W0.K.\#W:HGaPYJ
]7O3WQ,.@-e96Ka>]dF9;?=aM/BbZ:4AH;ZbdJ2AI-.>=B:Pa/4ba<OYYYg28GG&
,U0Z3K&B@]6Z83B=eL#d//FKbA9(9>7\XB[F(04)(+gAdg&)15PL(9K07Mae=G,B
5R_3\JDCY]@LF44VYRNUM/?4<LHF@-J_L&#8Ibc;JQ_cOeL34??g#f7-18[ZR\&F
c,H()2H;3Ed7J#;)@1)/bX[.7.5=?W=#eXP5N<g=(/3^MZV[>UYc\P(?MgFWM&^2
PE:K\66LYDTX<Kbg126gD=aUE5X&Ve#U+2ZN1:.fZEJd4g/41:)CNP6aOMNdT&f1
CA>=7R(dJ@G6&L\M.d;>b3?\eIN8F1dMH6VIAI8We)YY2H^fOZXfK)W-62:,MZ94
^GSO=Ag;.b<PBU+(Q7S.4:DKgOR+O^R,ec]+gH;JN56I^@Ye&YWJaR#ZM:1>2,9O
3[5dN[FeO#A\D0+IP6f73],,aD-H]1ceAWRKVc>0_C.e&gHCF=LA67c1Gg40YQ[9
WE9@(8BUVK)e3V.EZ-@WP[Z]LTWPFC8)-L5K5T=P,H1_8QY9dA(1A.FSg&C&.4,^
AL4YC/QLW@e-^aEbR=KQOG\K.P_-a\UbJ@.\YG-RZPATT>,feL^)^>L4</AeDF\g
g6?&;KH2c]85bA650E,D[Hee>-e@#??,;H)\bdG;a?(JP#@f?bWN9XYE@-c<UD_1
\@:OTCAPa=M5Fe?QXW+W6SUf^d2\eJWOcd\O\_-<a9M:gH2FPH0>JK,25JFI4];G
^&?IT/RaP0F.Z]g52,2D/Z4YMLg9(-1WKE=N<#XP7Sc>X8SC3B&X,=Pf1]MQFPQ+
]EJINTc&6.ILP@N/+=C>8b-;f84L<)bD<W@f>6RCZDB4PL=+Y@N+L-A1R;/JQ)UY
L,OPN0gM][R2\AF\SF5Ud5U[&CJTN^01UV:(b/f4=g]11\:_a?2EQ3gf&^3,>H.T
fQ;FBc<UZ-3>9FIK^P0YV?>O1#<-)D[7DUE5?(=D3I6PY5UJERGe2dAQ.JU8_S<N
3cZ3T1\9].=83QScF>QXOcX(&S6-02_7a,6_W_/E\YW;.I).?7<dR&f+EUId0EZ#
39TdC<8X-39C<^;:g=Qe:8Y7\3I?DU_/,g5,#/[DNCI,8))HJ&,XMZ9BE\cOFES+
4_AM<3b[9<acHQYH^Aa=:CD,8ZFOQ6+/?;NVg@\39>12IJa#FWdcZ>[&3+D:KXJM
]bB,d(EPXgbI[6:Z56BA\ad3N=bg,I&;dG^Sf@^WR_SCPL2-:1?7E09/YZD4X6]B
aB1\^C)7O67V987K@I@,d_VPZBG-=7@V\-dJN,T8dTR+6eB4H5feP]fZ1SQH7^Dg
,5GT5B^^2Y5TB9.U<H97-cQXa#>6/;g=G2FJFH+,3W,9;]R&78Y?b?A1;c(O>TAZ
dK]Hb07V_9]/8B..RM(<^UII[H)7Ug)P3BMSFfJ3f7\;A-FT)H()Y]6E573R7E;>
ec.fK8OP>17QI7b7S,JH9)80ccBM#\8WWfVJ)QTfNEdOaR2<4)OZ;-1K\R3(-AW4
Z7BX<\PEIM)&SH]ZP(>c:8V=3)8ffb+C7]b>-(SB^B/7@\-4/ZVI6b<a0e\F:UNW
b?fXcD+bAH4B90>MK:e4(gE6[4[c=AW@LK_DT.FEb47_<:g^FK[648>(,N#_[R8a
4@Uf7^KV<T9UFVCL:((6_&L,K#WD[:V(=IZ\T_+dA3JafHARCQ+2gE<DHGBKSZ[7
Re0E]U>N>:9I[04LG=:Q4H/+g=-FCFJ)I[H&]\@BK^OURHMA\AB:QX)47EX6<ELG
3#O=/EYA^O14M\?,CTUX4V#^-+,V,gJ>NE(Wc_DeHHSdRPHM]H-:G)g66gP4^FI2
[.JKf<3dOZ-1GF+2?\P/#:L[1I3:J<AcK)/dKB,=YCNS:5c\_XIbM-/)Be?ZfF2N
I+8\+LNZ&753Y?W8@d[/cVTR&&E5QfW,MQIFFAc]5DTGK@af9FJM.S64S[fZE/Y1
Y,/GVB/1K:BK]\RYGY^QM&LI]>BXEI_HAL\;=^c^1,6BZ1#S]>MLJc<XJ&((=U<)
J>D(BOZ-E2E1>PU9&C?1[f-]d4(#^D]3AZ&?;_W+1)YSV&5(^d]@J-DVR]gZGMB[
3X1Aa2BW8&f@<IgM8;XVNCUVa\WK=ZXfN.Oc[L#0aOgN\H8XQW.6_[CJ]31_(L/g
&81#(=dOeQ2>)QGVX^+&&JZR52GEf-L&I3+VJ[R=e:>4RSJ5T#PMD0I&QeKDLR;P
-^-=;HV^:>d?BINZ#W7T3F=,JRO:8F]EKdBf4@QDdVf,M,3-cYNC??Ze>XCa_)(-
BH3/;&E<4DM/(_b(JVPH)S15IA@QZCT44Vbd6#Uc3Q^Oe+bbOQ(8Ged8>LC\UG(-
.4X<U;8Y>Q8[G354MP+T-\&[=HJ&P8H45L;]EOVa?9/?SK:F+./dQf,B<&&@S.XK
IH+Me;O(=^@P6NIC[eWLK,2EGIR,(F[6)/F[eWA07X7eUSScaH-7c.e7>.G,+SU1
aaSN<cgH_/cS6A4RVaeVW3&@V3K.M<ISTR&J)KFUN+]&FN>bG]gfRHU24D6d>PXP
]3_42+RY<0_[.3_N@D&(,fTT1,aNI[L9FC2g26P31[,&dcXBLe38ZO-bG=fC_ON5
)(c;:PXbfUQeReAL/JVEW/P+88O@>:^:C@L2G)9S.[YRENV-L;_1#MXbQ1@;=5,H
TdWCFgBF(/(W\>9N[#W++C#H1:aZI9YB+H0XM:)0cXB4Ad61TH1AR>(<_HW4O[=N
PWF3FC/\e>W_c]EM@]KSOY5,PXPOW(617[I;fEUR#8J5\I)_4I4PcG>f<[]_[HN+
MUK]U\bg..EJ-a)]=(gJ+HfZFJ9]Q^8#7/8bZZDcC7b>1cUVHaR^N^RF?]<_8aKQ
R/@>/#D>D13bcRL)PFCB44HcKR,,+6C1H]9eO>IH?.2=cF?LRYZ<KR8fW:,C;4cI
c#^cdI9?5<N8+FRA2Q8/&5Mc>,X1A:#GZDP(A1a7E;WPS)1+GQ?VDG41?g,6c&]T
C&JFLVA\:TDgA89D=L6?fS>WL&]eGD>6P+1H2/M0QceYgPV^PG+7d7GDU@eP7TDJ
3DdKcGF^(CL\(>MF#+__F^0M+-=,cC5M+TA6^e4&95@0V.,c-gJH2G#GTL,3+1Wf
5V^-2IGNLL3cVKNa1:b/gH]J.#AQQ=e?Zf8F86De+EcHTEf]&]L2bEWXIT]P]Z)#
?[BH&gL,MU:fdQS9DM@O1:9D^<4HdO-OX7\J-GU-b@VN#;22<M>DbDgB<T0OCd80
@bOL6;J[=g7T0Y@V(fJLXOY#:\,C>0d&6(?D#43XD_W@=AcYI48(=Q7@c94Sg?0R
?D4,R9KE&([A\4&GXNMcET;g+813e#J@N&MCK7.OEFY-XTD>C\Yd8EBTTg)1LKAf
N9MYVYJ19gJV#C1W_0&8W1\./7F2LLKR-+<;8L1ZM21\KFH1@7R,WC2>:I]HRbg9
88beL_)1T2>[)[FOS;695[fIB2JH42^^]FRP>NX:FJ3J,Y_V2Z(DcZ<Y;=1H6@M-
QAgbc@/-9M?/)Sc2[0M-X-PBW_U^8B@,K;L.c-O_<2gb@FSD[b)E5c@F-EZQXUa=
5I,C<679gM8aY5+=X].N:CFJdTNgXGJ_B288J:[E:QE&28?V/LK:@5[J3(L;d.;?
@O7@bDg&1;cd0_8R;0JHB-S/M31KF+E3Jc0[,PUOP:[=L[-]=]b#4U]b#CP;E3O+
+01g(/0HS^P:F<A9Q8fDZ(E]741gfC95?^^8U0_3J=UQ\;G8ONgM_Og3&+O4\(;0
LNFP3_^81&-286/)GJ_6-Og4dSP^X?T;a457K(V0STR;<Y_\#3<;4H]=D&?5^F4T
:1P7,C>>f<PZ9eYD3:g]f96LgC_RP/T_0W-XR@;CFSKY&((P6F:4\LHe=1HGY+K7
0:7CR/OKYVc>(A4-LeQ?R+C/N,X7aG][//H;<Na,,^<00_fc@O2>+f9Y#D_c)>bF
@(BVHfVCbPcU]T(DQ&bK^X,/.48WCeEK#BAI<S]NLg3F<^?=[./PMgaM&RAD3G8<
YAD8GP/VE-T\1fXA<A?bL&dA9-N(ZacgIM4)AbRCO1[F78@KN?MX&?>7]=Bdge/2
S-?^=Q#K]?)L)5WDYCgLfc[SgXbD8CcG_B&4R0)7DIX4_@TTW;_FQIaYa&KX?63L
NKW#4YSSZ;BZbD7[D)b<V@9a-6Z800>=d0?)1AQQd54\]^B&Fd]+XCIecXY(I[>D
Y6BN:(U>b);\ZaUR#/QEG;^1C&ZFcHZ>H[X\OQ0>>#MDOE/.0U6BE+G6OHB;XJ,B
P7_/RB6#U)2WVccH4=NW1_2^DSG7Y50&<J;dU<Y4VT;_?O(,cBdg/UVGRK03P7cI
-d@7ON5::VM,:[-86_K\D<P76>]DUNDba:6SX1/Q@&XS9b]0U]^,^?;(dcTa48R#
J55N2_V?&6(0I;=&\S.?e3aA_HPVH5S2F9e6AddVGXb1QcFBDADSLC^ZEO-RG@cU
5?B:gKgKcdG(K4XTdD0PdFKS2;_LRb9FF:??c3ZbLSJ-B,OAC\7bN[S@UJZFMX:V
.UM=?8QQB9YBd=-VE>1H>]f=I][;LO^J_RO.^>+,LW@\XV(;O,_+;YHIgV>d3+FJ
]d)K,[R]\WK2G_f&1L3W.bcMD&JU4Lg&WPT(A^YRfY0POBBSbfCQ<be4AN[A[4[V
XX_7H9\@Sbe=4;Le7E\W0N5>Gec(J_O<f5?^e3+7Q4;\WZ=-JFf]X[6&GNBFW<&2
9fRASN0M;)&>D[1V+<,Y5:<]c4>1.KT/SYb;8;_:AWF&[]D]A\0XPDTN]_]6D>O)
1KX0HbWDMQ-K@C3[TO9gT+,U?c9OM[@P)TUBY_4JRMTW2@8R]<DLK=Y=NA6+LU4,
-N>LQc+K0dF3f861UC@gSJVEMSgX,<3;6_+RT]^RKMb//EK??V:d7)J5a#ZD=015
>J@2@VQ,P-BeDR2CIN=^Tdc(Q=P.<#A60(47;#b^\Xe9aV#YS5,6be6c7AA8e=_,
7:&N-A/KMf9.L>La=?_gd17F?AcOL\8@3I)gAK_OXg\F?L0fMC]N2QddB@)N:G_M
6XQ;4E;[/KY8#,E?@c=MD:#ZcaN2<@.7J7=0-O@.[2\IBMSECfTee15[5ZCY735G
7O^IaLX;KLH6d/0+;[GgcC[?SW/PV6G8G+@YCXE-^:dPg.W2/HOgAD&H/9?[X8NZ
Ja@O(faQI0c+G9.+-[Z1CUcOZ=-+e)+<_\47,K\gQfN0HK@a,3#PaSgSQ0c;S#8I
&_#CU2.7D&WM.H&CDb(b9gPA5.[eQ4AdO.2Z4f_RS0LcF\b\>AXBU8L7E<WEF+>M
2F:38\#3H9f#YDR8-]:d&M3.O:g#KP0+@XX>V.8T^3X=UR:O#8AK_&-MZ/T]QUB_
YT,YQ6O<(X3e]GTgTTNUM1E71b+[^2^@B);R_fM9^(fce0GU@,^74N/(XJ26cb1E
[M=>4##-.DGf=#Td[,QL[E7H?7[(eU4CEU96F^XM^\ZEeP]3a.>be9Q46g:D->,K
P/Oa4+F&:THC;TT25ZY)U=-D=X:CE]c.SG.f6+?>-gUT=,8YT;-R_b>Qa\4bd6[I
HGV_8TSc\;eaC,]325:JQJW&[UKPfPL-IF[)=Q@L\#beP]F_H(:g^+Yc7+K+cZaf
)]\gW:Nc1N#JHOQ=0.&,NeIB,LN69f,-M]ZG-.2c:\(28BRA=bY#__HDa?NDP59J
&19=T8S<A>\/#d:(K#9Q\b[LVfSU>Fd/bR/]>V\;)MS\NRc/a6DcgPeGC2;U#5-R
V2d(::VCFY;HC,(],Lb,>EV^@:?XJ,fVJ?P5;F(V0XVV6)::AbR94])U;A7][7f2
^5;;Q,N;G=a0CO\43cY.I-D//AA>bbYZg:,MD[A/fFg.^3QHRD=7gKcPYb?[IP(1
C++[:U:+-,?<e5RZ4=R:2Hf>?&:g:J6YKDT^G2NW.[9G<B6WKA54#V0F6^>2DWQ>
@eAMebU87M?=TM^Q=Gbf>a#7,=\\DbM-P19c;+F>fPWWTN:VG68<2<.,g+.bTB3a
;0]4a)2&(S2E[CZRe:N@X>)E#D67LZV-4.fc9.K0XCF5c/AML34&SYV4f.,8M00Y
L4dK=+R95_AFKVUVOY9B5(Y>89\\)0[VV8XeN5MP7Y5J/>Zd4;=O]V4OH]46OQXU
W6B7UHPIO+bRe&<UAE=P^2;Q8(@#Z@F)^T7DdJ<YWC914GA.dGGPHM=.[<H7F0(O
(:(Q:J]T)3&HLJ(5C1@#B]:2#M>8_=J)Vb<FCK9MBfJ\O,3d5[d0fKB\Ia<QT\=^
262M7aU>b^=B_GV+Bd]3LfS[.-4c+df_V#;LeXK&W/>&@0&8ZLF^Y_JK.2f-HU9V
G_KA&YdE4J.?/L<D0TM8dA@LVFK2]V9bd()HC+62&3RQEM#0(KSVYGBP=EG>CH,1
L2;UD[O>0[?c/SES8R5fK/\b6&eM.-.g.(-(E)bE8cSU96R,03DZJ?KYNTH[f3\F
\CP1B0AECA:?_14P/;6c_/BEReHc0N2#@2dbI&c;RZJ<6]IGZY41JH-4^^R4N<M7
[I?M3=g#e@WS5E9,_[8:.)M-ZA32/=]LAQ1KLP=/Q8WO.SQe#G?),McJ;ND(PL#^
/P2M(\faGO=TV6eAaf?6,7g+(SO2@0WVER2@I[a:=K9S^;=C(4^g=-IN]6<^+g5R
EI.FbcfKQSF0E[,d)Q97<7cH,d<T^-3<)+_eU7GY0I]P3V(KW[S?aO2BZDdOG>U0
+A\R2a(6:4VBZ9HPFGZ&9)1V8L^96CVMR_V00IQ5_7g,??IH6<>Qd>JFI+OA8899
L9ONF?IESW?H:=+V-G+D4aV[73MJI(\89>:B0&R.2+7G81NAL)0eafGO7:D_&UPa
c7U5A6X8J-4JFb_XZf5>eLMY?V(g=MHFI+aN,TQ@C9J;)3W#bLb\4d?W4Zf=9GI.
<&2(]B&8JJAU)ZTFV#T/\P=C9.J3]5_G,dg,Z^B.d&-<HfQXf5?941ZEC>b1X,-:
74;7Nabd@TRPHOT/59Gde[N3Z60#aNFe0/KN6[GN2YVM9<CS6>GcT\4Me[^_>+6d
.6:I@F^G1)H>&\]+,@b?YAd=ZII2(g&8QOC(g<F_1/^B=#NZT/(K@H3\CT9?QcE[
C>P&g]AD4=7/^\]X?S?96O,O,](&eV[NK#cX;@),d=]e[M81X+fUP1C6F(EcW<5]
3YJ(@,?QY\bG9<8c9@5#>?D/^Ya1Cb25O)5e,)^NRK\Z,SdEg7.X&e-J#a?BXO]C
E?^\DYD#2INII?0@E;BMYIgUacEH;WQ.&G;&IT-bJIc.,_]K=LO(D1E)H^</,),2
K,TO2cH)WZ_f:A&Za^=WPf^e3&cYF\#?(:BFU\f?7IS,@2&1=4@O71YK6Y)<XB8E
Uc=WW-D69)>BO#T[6ND:7dSA4V>BS,JRZ#fU?4>#OKFX=,F15c>cNP56?,+U7P^\
0.G\C>0UC^LeP+;F:S0eB#PV1=\]f?A^>PGEASE-1W)g;^]^/:<A68fTBcHP6NcK
R67dJE1WOeP.8VKYe3N:c>+G\\H_^@GR9)gN:W3.Qd;=O)@d<1Y[EXH<A;X1:;7#
S54^:&CDJeG016:Y3e/P,;48KB+++aVC2FMfCOS;+3OdW+HPN1F8/?;)g1HLXDM?
JGNUURR>P2b?WTRED]HCSeN:24a^7bX:(LV-b?Y1QA]ce1gN:?a0E;W(3)d0):IA
M/,NB+O0D>L=V,f>,&c6TKQf^IEI.Seg:[BJe-MK]LMa5PFIKI3B=W@PR.=@)Z34
8f5R2XP5@aE+[6GD3O?_5Z(P&BT1EUY;[gA]J9Q.VPWfD_cTI=<ZC8/KHL?8[X>(
9SP-bQZ;4Z.UT>KX_D:FF0^d.b3.93B2eM,4HEA3(P;a6([Z>)O?(-+]a,0Td+V8
1J_@=;5P(gLZ23L;]UWJN-L4G-+^V/95_3:ET/+3[\^P-TK9:bJDWR1+C4&dSD]6
LTJA]-R<WN.(T,UIJ7<\@4#g3(R7UF\_eL4QB+(6)dde)F6S5XA:(6+2ZIPGV7.Q
Z0N#@D21f.gf<CJ#5e^/U<<IBSO;VS:(ZI,3ZL^;A2///2M5\L_Z\?(;E6<\;SRA
g)MU&H,D0RDV,N:a]^&M@A:91QH#^QUKN&M#Kd)85FG::\_a8IBLfcWHK1KcW]T[
KA&CXC,8>-@7I[_YQPSN=f\#f:1,Yg^]4O#PDIg8A#+IYOd&Cf4B44PY84FMM\DB
8MYE=cRO/ag^<OEH[_TVY<\XUDe25O+61Y.][dRT>MW,AU@D?LOeM?Ea_D1GG9I,
(UH2g0L7/G.F]DH@?JY9@9BD_R,dbH(/R0a[6YL9c3Adceg@S\Vb[VF>X169_R2&
4];;M9F4A,@S2F@BeOCV6ONM;J&f(?C5.EV23P=+915J=<<Q42YMV,6^LGN?U_L>
:V01PUa<,OYFT\5HVCH+GGSW2=<8RS3R+J:5bKd&,@eWTQ1]b?:9GS]NY9f8&D@X
>3A@WSL/M>@=.FF+(Z.1#LJ8e&<(/,VE=R/c2#?JKCP.7?beFE0SX0^XOacS27O#
SK7S0.;#>X]5-^RZ.1a@TaG<#PO_DeHK]c+(#0Ff?T&N^8a3aEK4@f6#>D=fd>:B
^2K#?#AO/4dQV\WRY5H+e7446c(^QVVJb488bOBC/XCbVW1R(/DI_;1G8Rg07RU@
1fT1X.KZGcg=K<7\9=S22\75(XN_/f[662R<cDc?]QEgc>CGQN5gJ6@H\gcIT;\P
H=+VaH;.>2Dg3gY?=^c?:@7[WI5@bT.A+[Jc^baI]&(-P-?@77S1#UZ7&;B_3SP-
R8\6+63RKL]Q1-3=8^GGcda=\A&AO85cU7D:<940c>f?/NB3((34;8g-:VQQKNOU
HaWc@THM754<Nf;?)aYWKCIJ]eQS_PIeIXFdMR=4Zd3=fGVc@HN2N>b);N1O1(T1
<d/:1X0&A>?&^dO8g(g&@GAU2FcA#=BeX5Y05HJI&OeBaU,V)Z@UVec7gNK/7SX#
OGSeV09+B]6D)b-G@#E4cQIKUX.MO&^>3?SR/P)H\eaPX0aZD9\#[QCG,HX0HV53
6B:)Qa\54TBgODKXK_?C46SO;M?VME/dTJK>QP:565>Q@b5(\Kd2<>6_F<FN[fW?
ag&8FH@c=5;/:gU84XK;#@JDb_/>bFd7KB#96&__A182:\M2KcH#G:f:U2b7.92-
3PAY:X.4HLZS+0gA8S,H11d]SeO^EZT2_V+MbPeW:d(,O13I#SQ&#JN1XSS8N)ZO
<C>N:)L(YOOf504JJR2VN=d:NaB69-HPP)DK]WD5]8>=A^D(VWbI9U:C-#BGKS&@
;<gLI58cIHL+TVMN_7;bUcBD3HD(TXA[H&Y]AIIb<WH\&7;1N,V3>T9EP//AI;5^
Ca(AWID#37KTJYG8@/UYaZcJ,G\PX[I>++&aIN&5R>#gLO,1E)0S?-N6^,W,cLDB
/MD7B(7H>31L^ZTIU50S0^;1VMH3NR\2<)/IDT9F+E_?)R?(75f,3[GE2AX7E5;E
=5Qb[^3+D[E9Y8YUa5(@Ud_^/:->:bW9>M2:TYD;#OC?C<?N8RQafeOW>@KFCNHO
SVO3P>&Z<)/?[eE60_+#^MT98JH:(:OP09\Q4d2b<2PD.SAD:K]2AD[de6P;L]^Y
^\?]Oa;92B](7CTWb)81c-69EUJY/^bM7D<M0Uc9VUK]G&,HHe1geUMV1.+/-aC0
eRc@CG.MdF@M2eAHX@=bKJCP0LX+C[f@L4I]H5J7K63.J-gcdfS6S:7-0CQG_@H3
](HK[fcA4:AL#-[\B4S,;c@;#-3\]B5ObfNK&A\@MY0QB^Ud/.]0J[dZ3FD&I(2Y
0^3=4Ib(Ne7_4?_^[K.+.>:4:RI-.g+TG--4SL9C8:cfe^fO3d,<a6V6)L)M^:3(
a3:7PfVECG4:<Xb^f_/,C5_7G:.XZ^c/M9SPOI0)+(cI]+&C_eBDR[XN=7GH?#>5
#JdH[+6ZO9UI:9B<J5Oc.OX#FBZGK;>dQa^CYYQCVad#&ReKB</W>[N.YS+gUD42
7UOVC4)@(8^<C@S5Y-SEJ8^[/VAA;L>gO3GL8\OCUKC8N^b]K_DT@KN4OEZVMUAY
CX]I9)M8JM&WURD\FWd8]Z:KLb8-V=LQH,89YAWD&4(H3LD3g,Ueaf4;.g8SK/^2
(5NDcedBP;0S=J:&7RTUJXd]a4Y6\Y-59^#6O=-S_Vb^DY#:F3#U,O__2g(R/).:
FQ<NB[R/VU:ASGe.A+@(09.WQcQIf9Y8WB@Q\&__8SJ&R+R)7ZC\dN(\5ZXBI:Of
/6?:8[>MWbIQ(D._I3H\W==H7T.^^?R^&.ac>L,\XJJ[9F_V28<L0S.]W)_WH<^,
0E6#.Q_U:WG6FXY/P2B6]7URL86Q30W8[T[8a;BL<W)KI^QP1M36eJD1JUFN(\>W
fYF]cDQ\D=^b#Na)P3X>Z\<,#=UD&cXNOfV)--&D#?QWO&d;a2..C^V[7#V1PZgf
7Wg-P/HggT\Gf:Y6bDc=<^M.J>Q6(/5A3]d?fR]68,d_-IcQc/\M\WCMNZd]bI_Y
#+-.23459)IE5CB,6dG4HLB3RV&D>BYNB,;&FaL#W\T[>QT(^2S4K-&FYPNCTdcW
+)4F)BSgD)G1g<RWBQ/<:f(:?:eC6(A7X^K=0LNML8Q&:FXe^Y^f,Y9(2?5P;K(d
0[?69a9(>18^J=1;a)Jf)aGDSQCO>E;PHT\(O&G#CHJD9^+V1HM-KFP\ZSU)YD;9
,:.NV4YU+f<f>.[I]SB<_WTe86FT(^KPF+?e:9/2U;.DLN?P,]a4X-&;I7W_EHeA
4g/Y4]5>597]KOD:fY#YT,^Gf\3JOa=/2J^a^P>c^1ZYb79UL@LVE[XdC3aUZ;L0
+14-<CEK016UUSHP2)BNL@g\:ALc.[XK(6P:H^N<ALKX-NQJ4XK-GFfP2LTQQ=<D
4WIZFUA?T0+4Na+dOFWd;DAUR<KJ@#6OS0a2LUZ]G[+c<5cL_M2OBHO5:1D=dQG?
MF1bF^>KKD1/50?W-I/R8FWT>8:^6\&,FA2Q1-840L=B;+M,#)d_@CL^87T1#9-=
J0E[?-gN;NS3LY6T66dAb&1NW,HTAD7e<T8@(3g=\[:J4+7=a5O2g(Td_:>8/O4K
?Ag1=3YX,SF:7Y?YLd9&LabSP([&/LXG-A#:>RFg0=?H:0>OM+HCC&XX3B.gG;f5
?R[fK\_R;6&]3Md[e&8Y_E=5G1/L>4;eM#ET9U<CgSHPWJ.R8Ide5K+VW@b+U71;
aV.A\<Y@Ae,2:IG7B[E5#=C>(B)M-KG[6XSbLW9c^@UJO3,;=Y-E&-_WgFZ-0b[7
8_NJL4/\J-WUe.M-b]MaJ1HMSI>0)KHRMRO9?\F&:(VOHG1>.<ESVbccUE^:;1NE
DU35V=P]U8^aQAE@DJV-^b+9K0?cZVJUMg[gZT0R@:QIS1G#^J5HIJ#O&6#S3:(<
MY\f^ba#EdZHeI>2+@Hd9>fb7??264]Yb#+?6bJ3_-(]C?RIH5LQM,[d14aHO@SE
/O(OJGXIDUfP-C[X\C+3N)E,E_gQY.N?B-ERK/X-KG#<BF9dJG]c1R?a:SN3HU/3
d/ccL^SgFXC65@-+^GYN;9\).KFc\3GE4e@O)/;0,+J#RQL&dZLUILfc?Z&3#]0a
8S6cL@G##S2d96J7C:_;,dc3_^1\.6BAL\ERd8X?RCdE^P82[3eLfM:8E4Ea0,8J
g<+#8XLHOJ:W@0=HIURH#0Ya56M=Q5+aZJG/66PQ^;J41c]CLgG]FAI^[45g/S]?
<\SC@T^[^90L5;YHX7^R<V1e(<a-1OSTDQ8R7_\[V0YgW,6&I:4,_Oc4\7Ud+ZP=
,Oa=MHOES(7Zb[Z,7&W=(609Rd--L;;c+5<ZF6]HN^@^\d0/<4N/A)ZDYOG&H=>@
5_6G=E_BN<^bNC+b5[N6IX1f5/4]FP&O:THga@H@@GM2/(65JEc4IY-C&0#W)1M4
M+L,,f@eaF9K#bG>5gfM64FZKJVgfE43f>d7Q9f^6gF0>8RF0_CO/N.;M72f]I_W
d_bA@3[^34fJBb40RSOV@;8d.K^G21I<B#4AZUDb+,U1X-@SRe8IRcKP7LXQa47J
dXOPcJ0B0aU#T_@;e,<FgFgMe>QN5458@@3FJ@\@7<#LNB6[PdH3JWC9Ta3EMeC8
5;0>C2FI,5[R#UM8QN]\>&W)>49088E<PI<(eJd?9[XD6S(dI7,d\,<S.ZO2A@0?
C.;>56+5>?^Xf\6;@CXaG^WU>dV]-_>45OHg#G,J<[7CU<gH1NQM@,4KSF07U2-W
H8c1^<LS<+gI)5/LbQ_^W(F^,<d>DVOL(>B>S/e97<6Z1B._MXUa=cF)6.,5:3XZ
YP]CO^,/(LM?#>EY2>L)_.IN;ENJ9WF_.8PaNgO)dY4&a-f+]9PcE:T@JaU(\HN<
1_?>fO0;P<CX0<30Xec,(4@WX]&;VS<J[-cF^()E=.2AQ[,NVB#bFPPMISDM,VJ[
1RZG>cOeG+\+]=5TH4BRdF.T+-e&IHV]NZ@[+EQV5G0G](X]T2HYN]3=_5[?ADLZ
QS4X42UXB];;6DKU\&X0>ZgAD;ULaUeX3eN0E@@::9,b?6\2<SX\NKeaKc\8_(\L
0+9a&L&5C;[fXQKB>PO[)0Hb0fFZUa3)-:O-Af/.-EQ+Z6c70Q@M6RE8?-N4QT3M
MN;cWG#;F/)fWYaVJ2Sc/>R=1,]VH(/1(N5NW,EOWK]XO4;82QON75bN[)(/VbC<
gFKLWKO4T5D?+f32.TLC</g[3[Y?R<.=^MOPVQ/3ZAg=QT37#1EORYT]R1J8&bf)
.IK)9IR?Y46_^B-SNSGDCT-N=<a.G,96[\ZMHcB4XERLN.Z&DX>E^^6T[;^Zg&66
V5S>/M/D.DAARLfMJ_@P27HJA/=DIGfQ+0L,K-bX0#&JH50DRJ-9\N=UM0R&_c&T
]O9CBA#TR(#)^:cM]G]<cJGf:V,:W(a#0N)UeZ-]S?K;2WOF7^.HYWBfFA9V+P.P
AHBQ^:_.1W2R:QM+FF)9JFb(AJ+SC-13e+&TD2OPT^/ISK135VD.@IeU9ZAN>f:W
G1&/MA9D&.d.RA6eC8&H20)#7I1Ne)^3H+L\>cZWESSIZ;BL2=9VK>(#^N.K2:08
:.edR_9/5<UMXdK4?7eSU>c<E+IGU27gP36++bSV]A=/N1F;,af:SIgZ##:D7FRN
&Q+XEZ.NdO;YHKUGF=G;P===7bX2:1RXVD);Y2/<5KA&_-P3<BJFbbY@:F_VSGFI
Q<>1eZT_2RMT8f_e=aE_X102ZaC4(_0?G9,)5+1\T/;00R3(a7?>EK&L]MS(=2?-
^QS]F6Ug5MW_71D70O?<O1C-N\&8+&+8TWG]9Sa2+R[b70T)ZND+:Tg_:DE[\-1D
[aT@bEWXKGZ_PVeK5>JEX7HB_Ff7IY(D<UcX=]0VKJd_PIBZ0XG7U@bZKX9K(Sd5
?J5#7A7\(4/]J>5&MVXOL>cB2\2N_B,5dTLH&-e4aSPZc/FN/JX@/S9Bg;-?I6\F
>1\g6KVV-d+RcLJ-XZMP[8V8HO&E?3D;?73QZ]._7:aU6B)^1&a]03gcV:_b(bPM
E548RWc=_BVO+URBA.+(=7RSAP?b5S\_Dg;ZQV#5FZH+G+K-(5bcI>F2TaWD7+NL
-&2A>9-KdZD@Ae;Og3;?OPR85H=71^J^d(=C^Jd+e+J\>Fb0XJ^GFJd8N8I9_#-Z
NDAMJ(Cc7Qaf>I&Dg+^5A;RP@UgEYNbOR.+#9RCSJ6dP4+4=QGb4K<98&7OALIb(
&VKK9W(9;,8:F-G[aWKeS3>FbX.gcgb/eR#,T(gGH-67dV;0bg/+9cT/CcU2OGW(
dP(;^>d?KG)G^N6KI_\7+E+T8:QR-7G-+g\>-BAf_?b7\G7E^.]I5d)G2Z?fML7Y
2:8XV8VXEL#P<B,cdQH<HN[aa2gA(H5,XJ?HQL/>4PUAVM?@0F9QaT\0T-(Y]]D4
S(<>,G=2ZNe5.(eD8+LB=e-/B=cRa^[&:=OE=+UTW9RD]gBPIV&6LCVJ3#Cb>5Y0
)^YF/b>N@9,MSPAFLPRR<85c82ea<KL\Y31+A]4/e.JQ]dbd7P>0cCCVIb.]YMDR
K:7cU\IJ)gaF0JEU:#?B]6:XH9NGfRF]I)NE0>NL:2W3+(e3RQ4R4=HFO6^#2g/g
c^Z,.E5=AZUHW9R?a?]W8bY5\\3DG:G8T2:M^@]T2=4(K&\&L-7dVSHQ3P\LH.P/
,TH(NT\X-<aNUf&V]S0YC=R31NT?>N)02ICcJH<K\#U:fCG?>c>?Vf)09K/@HA>N
7/@WPX^@X>DNFVZ;^NSY=cfT+82J1.?eBf0@V]GMa5?0c-X6>g,^]eP.L778H&Z(
&:H-CL]7aP^5@P-EdR(c,4C]\8MMUQ#BEQ3UJ?#K\@M8KZ-NIaZ\.\S^57I,ZV&D
1(8@23/<U?\SVJb^)Q_DDeL#gBP_XV.C2:7051^Q=[c,:1&1>,17[&;G?AdRZHcE
3MDXP&9,6VX+KA<6^fAa<RXTWFM[5?BEK)BG<[4.eJ].644ZYFW5f#_4,f3HT/#T
Q4a/Bg8(6OSA>(T_d]X)5dWbP3YXM=(AS61.W\T:;&Mb\W+[K0&)-d-&P:6@[#IL
8S_dANZcXG24dJSEG.D_T>cU?dc.:+SgTPf>I3P3+U9JLA.=5:>[_6YV5/-NU.B;
6G7BO(e1-32Y7#RecSTAAU;S]8TKK[-8e0UAV?D\aZ^b[SXKPd6D&aFaOK;I^e>d
<]Q+>:,6+L(Z4Z=^62PM(]>GS+RQa,QcY/<J7BJK1I>L?2;][W@NKde8/6Eb^51>
E)T^((@P,?0QGPMAc^V>6?#XJO48?)E6?LTgP3b]KcWN,<GNNUUD:>c01Aa8V?f)
;<LE&Z.D69cJ-+W&=?.^Z&fUW,=KUA+B=,8K7I9fI:_CD>1H1/)95_8EdL+JD?^b
+#J,_/Ld9=-S;\3b)IHB(g@+K]WE3>#N>(f:PK\73Z9K>@aMG>TD(gI(\_3[bM3S
EbCad41N5E6QEHf20Xg,-[RZ/ccG-JE6]g#U]]O=SD\SQ6c@),BKZ73Dc:dE[.D&
@9CDcf:H@KVD9--3ZC[2^-Ad\:b76_5\M:F3IQ4&I.5E.Mc^)GAE^@<fNS7[L4?A
M:]V6US+:aV_-&QTF.;Of[,0V3L,PAV6O-)9Wd?M>)\,N^;/C97;Q@5#T5.bf]<]
&QT-GQ&DR:YgE]J?W2_F,MFI,c5W]GEBIZ#,aNd]\+JDNH:Ga),A>\Mc9V=WbH,U
1[C0RW>@Kf)fVET1IgP04^OX7V_V>8,SHHMW>J-=O3NYY#^CDG;1VD(1VaH>-96)
ZfV7P<Y3@,9E2NCZ3<J]1X7edQfCW@,1@IE[fGFB?.gfQHRG[D1K)0VScA9ddeH5
P.N8>#1_4adc<JQ.4baJMG(a.9&YY/dBQ.\.E&HeE(F1F+0>PZb(Ne\Z)DI;63<Q
#PeBXWZ5Y]EI:WH8]O0(/OI>D-;9HXQ=GEK\0#ZRC/DgTeFU.3<-ZM]Fa]E4XKC7
=K;T+^2La?RDJgQ(c\M^P>\<P8E,6J8F:_??\:S)f:81TK#SW#1ZJ.J<<ACdFB?\
DV,^_=4g.1?9IXRO&abR667M:eR@OK]4]BT4#gRaG\UK,/0=/1&O#&QQS3.#3CJ0
<+L?TcP<3)_3ULOMTe1][;0aTV7)fYJ5BD.DFM-9f3@R5;1GO_eLFO2^C>>^f/Ee
IRL>G#;GL:@cdbC&I\NNLc^T/32E?SSR>1Y92a=Y>:G[W]?LM4CDBeKc?4GK4J+<
+N4_W\>Y29a9^?WAK2R?5\>HS]SNCM=\Q&dC5.g;Z0#_3D:1g0<@:Y7,1R@;20<7
ID/T3;8CO/+<O@f(9X:/>KO@8+#@c@18<b?[&WAGWADU;AT0Ad.5A?Hc#>Q\1^R@
CbSW5:_3O3Dcb&B4VV&8)X=/36:__(\8YbDOCa?c-Zb>2ZPa6UUM@RaFdV69(^(S
Hc[VZ.M0/d48T([S>\C]&9Q<>^2ZeV>7UCV];0]^g^ETXg]H19-TSTSV/J1cDK=c
1KSe&F@A\TJ_P.P0P_Qb_;C<UB94=Q9L<;RRZ7KUBLI&6cYMJafH+;fb[O3>UZAg
35^##AB37]4A(&cF0&CAJQ3X;bcbVF8,#F+T)-R7M/(38@#+;M@dMV^e)N62?52c
W+0C),@MA3cDBI@#@&^^,2VHA&15Y?=/P5H7:#X_D+X@B;W>(4S=2HS-ESd[<4_B
Z-?Y#S8Q\A+FWYfFOG>K7Ic@W^]/.PCFN_:>8\+;E\dQV1e\3&Gg&99Y^VLcA/Ud
[O._.8,I0^OXZB5+Ig-(;<ZC+Tc.936Gdc_@@FUH>U56HV?3LV[0]GIe5CZUT+\7
EDbaL-GI6Y\@S4D##746F.Q[=\GZ0-L2VLfN<7=10Pde7&Q]71?GRUZ8Q8dDZ0&E
E:U;Ld1\:bM;>C0U(A^6#+#<We770f-+/.TEI8&VeD\M4?fe=MJL=K/8gDSMgQ-;
/YJ;-;N_R0SaT^J9\X8;T<KW;()D?CS:3?)T1e]d5=Z,E;6^91ZR?1F8@JA[:ACB
>6UDZQ?Q<GUd[D;F/T5BCdc_d7E?GH)_:JDAP3-bWd;a:<XZ+.I<<VC:E?#O_.AR
OC6TAKgc&Rd)bBF[e\PNgcZF_3LCbZ.#4L?gY;HBaK;YA7W#2QZ=-+e\SUZ\ce+C
<4J<?UJ\-[:;-F@5ZNaU\26=]dcg)T.29fZ0f^,bbgLZUgB^BRHa3E?UFWHN;CO]
eNY_g+QbY<O3_MW7J^gJ^N1>LKRTZ1:OE@4?7HKO5[[AMGf-C]MR:F8M[4R^&YH^
9:CdZGf(9O#7CG>D>/@@d-eCB]V2X6eYM9[RG_Ub^>W/(c^YH8\e:a6@4IS>9:V-
6A9H-(_<:0RP059+W\#<0,Z]e0L_)])BA8648>e?J&d,ZgN]?8):&]AP72)Q]eJ&
/YJ#_[E4-O1Y4?.G#/5#DUAGT:^a-I#HVW#e2S]09.<5^Y_=Y7(D(ZFf=?dOQ8M0
A.e-e)F5D85ZBBPXDB9D6J0XMQ3aX,1g=La1[4Ue8c<+RMY+0e\]]9S(8Bg\#PPH
[NSLNc@@K)B<\6[DJRb1c2#HN,972gf>(L[^--\dRg\6Y?J2/Y;0NH]JYg=LCQEM
#V=JLD)X-JaI45_0gNME(XD5FCR(E2LWdgITZAH_^_L_Jed87M/RY1EKCEUOddfQ
\5@GI],Vd\B?4Z_L#.LQYGO:Ka:<^)KGX^OZCDg]]6\FYS^Z(VgL;)]Kd3IH#LQF
]BM6K/Q2EOJW:>&d+X\1K#4ZR2CRJ)M/;[[L,U)R/WXH2BPSHNd0?5-JWK7R9<@Q
\:Df<0,T=aa=[8c2_.HTN@B@S@EF)_aC:,0XR>cW_AV+NA6F5>_Y[@JMVZEa:G7a
.2g0R&Kg:8<Of&9K]&S>0PMV)8.07D4S-8:aA[C3fBc?,XXK/GPA/bD)DQEDQ?6^
S#Z0bHfNde+Q)#P,Kc2+\/0:N;87YPLAR\-@HJ7,9:IEd-PRE<405,M9E8+2R/9Y
>S^aII,M>V24@f8Q#JfC>-H6_]VTeVIL7&[1g/C+^0g+O4H3#0:]P3bL72NF&CXQ
Q##5&g<FFe.8(.IZP1LDG8S1C08^J,0KN7G5MMWIeW1=\FU(D:XD+I,<3(8]Bd[K
5(.=7U&^BNVH>DF:W5?4[>GS9OHSa;)>gbK_P1QG.Q7M6O?b1N)2/#E1&YM<3P?@
(a>=WG[5^Dfe+(9:^NUI(:#E;7S#-2OBP6fg4ME+X<>e)6<<;a=F[-KL],0I-IBd
>H-<JUKDS7_d2LecI3JGTZ=gD8&5X43B.GRQX-bQg4GO#<PaaL\4-gZaY<D+Xfe=
/X-dgY3:e>E<[]V^]#=R<gQEgA8H54XUQQGN<>5<XAgVA[MUNe1HN\):a/)_dB-\
gE2cJ/d.6a#^C2=U-60,CJ:S-Le=GIK-aSTd^+B?^C1Na9UeT](OA/N1W+4R=?dD
f>Y@MIA3.46/?fOMC-bAYA92Z?\cPbS+e-IWVX3J@cc^\(FdXU-?[TYDeR&0ES/W
S6LS@A.#gI,4Eb>=IeZAM6c@D5KD[f\B-^M+-e3CWKX:5B9R[X?(&f1>56beL[AH
I(R@[H7<X2.&G(/G<6+^C8_Lc+JK+gR8F>P5d=)3RB9@^,-NdOJDT(HLL(U1F,EL
3GJWF=c<..EJQNMYcJ^cFYAZR4U/#1JA7d;;Ue3X7>MdJLN;NK_e=g>URNV0PLY^
.&UC=;d]O6T63,1>QTbN>)ZbdZg3\gOP]@N6S+SRELZSVA(.;\W\S3Xe):]A3L12
I]>(QG0b6c9_AK[_AA^_@)\5,5#^cYLb)K_+0E(-5fVD:HeFD)W)NbU,A1LS+Q3R
JL:DOcS-f7V[b6M??gWG&f]M)+c2Jg:CORA];I^SUQ(:>PWH[,4B[W]f0Kf/0Q?W
fW_N=TYC\THR32#X30<?\433+Cd)\@-UV\^5\37=4=bIfT[U.R2^7fTOSNBGE^6e
V1.GUO9]66ZR=fBC#W>WHGcFW+SK-LMT=4@M3A^TTO+E8fD523]@?K+-,)/aF0:Y
\V4WcKfF<+^DTJa.7KOZTO9cCeM.ebA4V8^@TS);5)#UU.g1,Kf.[2)G-;UG1.<Y
ZXa>YYE:;#:?80=]<ZN.?BaL.D^G0NVJ5f;H&XJGI3IEL2B/8_4(8M/;227/G,1L
(2CGa5/_3/\dfAA@Q+:KNe7<[/TGZb&g6],KC,L/]G1KKR/2Y,YW14]Afb]7Y_,.
NfM(6SY3RZ\4<W[2KL9?-LSg2S3+YL.eN]N1XdUS&6N\5]#<B3T=#gC+<-)UeHMa
IUJWC;:d<N(2]I,O,GI>Wf))[K3P-cg:Z6CaGBg+C3U2bCVYL(Uc(WZBcUQ\)gZB
Eb9#ZR::KC1aLJd)cO@0TKZWI,WIX-3\1YVP+9R=2&,GY=@<A-O5G2LG):3)XY8Q
eQ3Mb;a#f<?dN]]=E.&/UAPd(,S:KMCCf<_c\aX[;F0CfBMR)T@E[V0\Q#U]b/0\
ZS5ON(\.U?Pf(=/421ZUCccA8@PO8I-3\H2.:F1>S]5D3&D5bH;)f)E.?H73E:X9
2g\b/?8M.X_P/6PgX9X([;J/F:;FBL-VWJOVA@O79Q#7Lf[Xc-1Se;RcM#MM^^IO
4@dW)e[]6fTLAggERG0TAE3Rc[d,=0SJ7cPTe=;5f\e4V):cL3T]@_O/Z_OO)FQP
PLS4<TK(^@,Og9;R&BI-0?/=X:Dg:N?CFJ7VWO5<,?]K=(U?,MT>8)4DB>H0\?1D
YLUKEHR<V[L&(WRU:1T_ZA17\@(^4&4VM))b&0;34666L+;L9G9P\\Pb9P-2,dB3
^CA86.GB=V)W(&N+G]1/QY>DB>CNXb^I?=Ne]0eeC#RUgQN=O9LgBagDR8>7XFQ>
;B2A<[\#Db68W3FYR)_H;:][[8I+bf_]G=(>T?^K>]DQ9Q_&A;]AELgcZ&b42@J:
#f:EP<G=@J^aC<\,;P8;TIIAIVZF]5TQAL.^FR<VIa-@bCET[?1O)?J+0e=+HO2Q
W#UIFI;34L5dKc.Yc<,I^?9X,D^;5,aRDa\#?=J&RHg4TY[F@<U3PTAB6/3cUC__
.RC-0P9Fa8Y:T31(&;I_O4L-OPa7==KSEgB15#bSF9F\499HBP:2E0RF.ZAY,6)7
6Y06=(\_IaB3#6[X<^2aK[b3fYK:NdJ1QAg[\DD3BGdg&[W;RXL_dC4V??d:AW3M
HOY3YLe\BIbaY,,QTcRZ904J6A<N7QZ4GRDb3ID/YcIF?;6G_[^-TXQDL\LTcBPU
U-C0A0B8Ef[BE96Ec5;M8ga&;CE/e=1[eIXeKJ^\gA:@OI)TbYN=a+P4Z,CM0Z?W
f7(T/9RR7]FdHFZ#]GVa?JX@>,X=QMV,1TTDIM+^@Zd:LAgcfbPKa\\;ACT],7T;
O@Xa03He3/Ha[b584=3gaVIWX5)O+LBgF[,ROaaY9@G&CNQ].b0@Hd+Hd;^+^2e]
NgB-=NdOdS^/[XNeKVI(<3=3V>OKM_R)7?;-IaBT4R;^/8M3GEA\7c60C#NJMF>-
g1cU685RT>b;9]>g(N[:O>NAN?,XBN;_P5QZ8CaO#7+FgS9_XVDFKQ0b=b62N?4a
W]\+Z,ag94R-eQP4;;>RM@+XF@?bDINFHA2()KQgG?98]J<#,HgcKR+[AbgGKT65
I6#-7=[a?<ACJHU^IgGC7E@1)PH=@NEP4VcY3@CNV0f([W5R)<V>ZLg@=8C9<RTV
CK/D;K^cL2.J(EC4?b-g+9\XUN^QZRO9+X(H\L:_^NC7L<eOW6]@._BX-A&5^X/S
5aAU,R8IAKDQ&2b78R/(O(7I[B.C2/6>PH^de.TbP602J5YA\?&?ccRO,1BPLeT9
G[,]f2ag7TKa.(IWg6e9Od.;[RPS1aH,<?68e4+[8RG4OIOU81WSM(]Z5+:;XY:E
VfOG-<VA-fgd5XY4.WP-K-g^U)\5/]2S5)G^QbX@fOFBI=NgL53]&\MZIQ9+OAC2
S4<7E;_1[O6&1JGX3dVL:7c@YG_]\aO@dT3JC=_RK=QPJALFPP+:Z-:>HOU?(X_c
3>S[UQ.T7B^OYP)8JXE:K/8^5P[e7U;_3_K50g>cC\3M=O28T8=A_cT61a10;SId
>8-WYX<[c8C6#[3WPa1#X)_Nc3JR)F)A6B]E+:@FSEPJ^YgB?[1Pf.KQI-/+-.<&
T\T0b#dEEEB?)?X5#g_3B;M_S8acQ+TO?C(A_HMR-I#1^fb&Y2Be2#^S-KB;\bB6
Z/JUEJ3eP5O1)RI_>8JPZ/d(_c,VZMed^E[aB6P;IgI[-e67+?5&3<OFGdL<B9#Z
/LN.(3T<0YbET,<]d4/KTc?2IMFg_7Q),L+9YRET0&I>_QQ8P1@0g__5.JL65FUW
JYb(TQa6e53;G8?:A9X4B2.gFT@-eRbA)5/<faFcBb7.AH[XFF28WXdU4.GC;&D#
E3:&+gd=-_7(\9T/9C:JCYQK38;BL&0+-aZ:]&.SEa2UK\_3OWab9?[4G?9Y7Q5J
>5T(>#YaAN)>V>T4FBUA<]/\8&S23TVIRQC_IM>Jc?&#3L_8;[VJ@cA/,KK,6Q0D
Ne@@(M#C#&XV0A&]L>F#T<&[B3fYX5&))Z_U+/44)NA,9KA-+OJ0HXGL\fS5eM3:
f>X]=W2.[-c>De]3-A[TLE2I.0L5,G7/cXJ<BfaU&2JI&_@<LC4Z76W?:@F6Ug9\
/OUR2+b4<S+D)X)+f.YAb.8):FTLFX?N,US#&6?HYC@/F8ZgId&C^IUM#,HW336T
KP6BF#cQTMYI\)U1DQgM7;AdA,ZKKJSFI1H#Q9ST^Pb2b1b#1W^-A0&e_f8KJ9?<
^/^M>@RI.)4cDFIC6^,T3^U5VYa/<KL\RIH4bZ-c?6CZ.K6O)B?MMOQ7YW@PF392
b0b#[>MZLeJE&b\V)bJL=80=OAE>A7.@)5Y+cfY5JYW[903O08ARA-PSQ:\K7E2?
?-]ZLI3Oc@G2CgW-36=fK0a^]DX#70U-:DDX3g&DdB\^#>;a)Z1]9>#/[]N(--Sg
^4S(HYO0(8)TTT8+e?:Y^YFF)(R<F3[;g=)ePV9@MMDJYS/=A/a_e4(RK(VCF1Rd
7<E7__eQ[cf9LCZ@d-)0<aB-GI5^26V#?3.I?a@#>O=\8RAWc68T@B-gXg:I:GdG
E/;KK;X=SJZ(M^31TQZP1>\gd2^:P,6]5&<E1gW=R;#G;XSZFHD3ROG^X2d;W694
<Z=VPbd6SVd=(J4_-4=Ff>>>SI.1LB&#T\QDDE4+_#F5.cSPS>PS-7<6XWdT-D6(
G2/a9e3889.H6FSG<S[Md2K9E>cJV\SD6N8^D;G.ZNRISR<BI:>Q;2@PR]AW07//
0XDcVQ/5EYZa@X?b1.:YE;8S@VDWA@U2;_eNMMVKNA+/))Z9Sf4261@:a]F(=L6G
,;\<KV4U&a@8R>9WHHP^++Z&^d\>_Z+[cAH<cX/cT^K<=Y.U)4g0SUg?f)+f:1EA
)76+.,d@H73<W[MM<O;Rc<0@:K)dfHT82a+]-?FF/0aePa8LF=]7DM@HW_0@[KIX
LDI(a3cX8>@:)IU)QR18,MOP[Q0#4D(F5@Me;_\K,3^_/\+DF.M_6<afRP./U:c^
]&>g(cF:e<J#SEU/W8+6RX&RcKMMOTC78=1=5_7aE_e?@:_5dcMC2)P(J<Bda\NH
,)NT/.;P_B[WK&=W)TMAH3-_A-EbK3UK&/0K6Db6Zec;>/J^U7aIJBK^:=\?<eH>
cCe2R[31XTf-O7H#BEW5JX=^CC]E20Yg)2KWNDL;Bf;TJX2PNQN\e/1210KXPKe#
+c3W>]&6MN3N=GaI:3?CD1N161BU/:)TQ(Na^+.?C/T@^U#7#e[WFY3GO]7F2g^(
c4YU#JNYNL3W]PQP-:ffTL=:4DG;3N,=b\bDHW@Q4T\L[_F)N&cH7D[:eS^@/)eg
VWgS,c<WM//ZU=TR_]8@-A7P\19^J.Q;FH@NSZ8<O1LIY69\0_7A//&gQ3X_B4Cd
K834YVUA1C^SZeI-:T@CC0L+2\=(Uc,8d_PX5G:)+9]QWcZADD&56?BN5SAVKCeC
OK;IFcL?I2+M/F&-+.Y3Dg3S]GL]G&]#8K&Yg?1g5VK(R7/A.DE-e3YYF4A/H>6+
DK?S,Q)bLDX@1VA^+I8<&b,SCNg:#:gWI9#8\dY1FgUY;QF-?)ZL#X,GA^VETUe;
F9X(RWM3@I8<d+0cR1)EKc4FWB7&S;CE^DX#cE<V[;:VXaBK#@A=Y1LS6;HH9/]#
?05)KB-e>9>fX9JXg7=:6e/JRM7RPQdC+@,cH,g8O;GWOZ?TdA,U7d^EF>(>AG#7
U?A47Y+G+ZN:JQO:^0#&=/;GeHD_;0]L5)II&,&A/>cEQ(EW1+2)54W5+Q&]<E@Y
>N.Y]a\WTBBD=^eJ?O]@<IOB[c5388^5WAI^+-=I.KGd;g&7J_ZL4GJ5=3c;3MSG
.,Zb;3@f7d)>[IH.Q7QK3cNe81)c9GVB+BdT<g_E]Q#8::6>7:?&VXGCfGF>_G+4
=_V=#_A\g<K6c=P,<;3_dH;=)+-H+c9fZBPK:PNaN/=:GPDAJIR;9+-=I@<+JXOE
P:FXg4,[:]A(1+Y)g9e8SZ=LM:a>?19f5_S^)ad>IE01U>QCATNN377,3U7,<I)L
9IGL4O2H5,g(2>^6DNCY=(/F[2E4YV=Q/Re7;@dSI&\2:\^0>U]ZOce.M)_8\7S#
7NW)^B9,bg1QC5E&B;c#IRNV5:C9a.D]<MT5ae)BdJL_b+2[L8gcO.8L4#,N,S^=
0)>-=(IZ,NHE@]c6OVGQO^_/aLI:QPPQ8Kd4<BM>Xd]WCXb_G8GRE6RYKU:[&E=C
AIa?;R,@S&H53^9gQ_DNR&KR>7d:eFHeO_=2181]9U);[)M38I)J0.PF->eN\>9D
G8gN\5BL5EcNOZCeM5(58A\f#_6Q[@K3J;ag-3bbK9I0PaC:1C2I&[Z]]#)4TbZO
>H:+3A5YEWI)L:I2,C[5+CC@XCKV::U@.9^JbOgO?W0;)):13>+]XZC#(;64KR<,
g(6,b:),YQJ>FBL&G=_PJCfPQ?(7b;A?N[]:EHY3QVe7&IOU^<IIRVebdJ4(I=Ff
<EaFEg7Va[AG<B3d1B<G^P4?-_<WY?KW77]OJ4H>S6?9)]K/K@LTG1]#0-/-D-:f
4P_cULJ.)L+G2O:-g@J4+8LP)#a<e7aQQW(gcX(aL7Ee5#4EeITP,&Q&?<D3XbWM
AWR\?e\D)_PR=)@,=WYR5FOYC)2<L2>AI)BDCL<SB&DX,9SKQN5?D^?7I0JNUa7Z
?7;#](R&9=?2))S?;&4YH;BR;-P^C<M1,=FX0@.,^:WICgF/\?,3)fN>:CE,EgI<
V2?UY/8Z8\X6^Q5T11VLFW#(F@/?dH=[_KIM)fDM3Pb\2J7NR6<D>Ye,#)5.<1\+
X2H9&(T9@_/NMWB(cT64e,I3C=fGB[EK<Z8f>48>)c(\JD845:fO6OfX&&K0eZ-D
bdc(+;YMgIFYAZb_B+M9_cH7L^=dRD2)Ze>OW6YSBCJ=dfa>eLa3&5[)gg1b)Q_+
b-4QQaV_XX.))(U-W;>Z4Q^DgF6)G24&&R@cM(#,V7DYG-Fe(6L-)<@I(;8fNU[9
/\WAd(0(?/B\W<O#PF[MFgV9<R5[>dE,:CZRe.K0J<ABS<)]Y00K7Q2GLN+V>_5A
9)OZXFP:7<Z+c1:(YFI#HQ5W/BUU([HZF0^&XPM(:3Z8;GEF(/-S0;G;aJaB;K<@
S0R3e/;2gA3^+e/WQZ82-XRX/YXR,/gU\#L@QV[d\QI+K=E](E(:3GeLa1+c[PAe
IN&g_)(?,YIAAK#HSZM3dCFLb1:Tb3#E9T5]Y9bEAf/@=-19@FIQ/HTeK.NUe]\7
B3cF1@HcZ.Q^SX1C+a:.)=VLGADdePJCGd4:DD2AWI98I8ZGJRKJTF/b);F?MN^2
=eRB6W6--8T?1e=7a^X-f(#-0J:#4>T7XUJf0@3:Ke/CL(1D)N<NF-e-YDW;He>K
P=E>)7/MIFaDPKMZNE.[OX7=_RNS]cO6GZf3g:BSNR&7=aYE?;#Ee)/YY4cS/XPX
AAZc)-[#2_5/9U(C-CCWH;KJ^f3eb5GP]Y5:R.OQ9<GUfXc\05Q??/X9aK>6Y&EM
]_R<_TCaPL[4)Zd?GB+D,9^@9=eDgOV@_e9eOPd?.K@G;Q.RJOQ;Kbg]C)[C&cVY
SJD+f>e\Fc\1F_Q>60YYY8fG&YBS?L6/8>@K(NIGLMQO]D#fYAe:,>A_UbT5VU[9
K:f]Rb2KXJ1E>&.-:3f\JZb.b@We9Pec&\XGabH;RB/HWFFS<1PKWa1,+]^LeLFQ
^T?@?A2>)-aXNYEK1R/-5;I=E/F1,47?5J0I)>aBbMa7L(M2AHUJZ;VOD0Q;Qa7>
A(bV<2?BCDLOSa\:eJ_)U2X/XMc:bN&\H9],gg39)[RC-W,3HD5H,G=?>[5DL6<I
):GQZM+W\-Z-DY#8?)(eJ#6#U+F#ccdW#Z#bA]?;:?<+D;CFff-1?M[f-8[02gNY
YDGUNa.,dQ2De/;e1&eW)AM=U=64GVaMSIU2[ZL6RW:WfB.Z>BKHK@Q12gW^CT1V
gG@J7^[F5EEdaJJ?+.?T?]KWf)FDEbEG:[KQSHcG-:7,(9W.A;07XdcU?3Ta,OcB
N1AT>::=8J_?;:H):YGG@I+A5cb5d/H]=_,0T0(PK.?c-]C;Sa:.@.#1aMLWVI9M
^U8B;=ZN_fP(/.TZGRaI,U5@+3^e,73[0]a22N2)PB3?;=6V05/_J9SY;T3;ZfR1
c_)LVc3S=DbVY7GeKCAfD4DZ2/3W;eIdg4+GD+g<1=O##_XRD>>:)[>,A&59V[8E
6Y;93?0(Z1fT#;JdQ76M5aH#8.+G0E8d7E;.1T<1\1db2FL]A?]3WXf8@47D_eN:
1BE0OEF_UgBfF-:/1CTc26-N4W,X@C_F7GaDG/28>Z2@+X_GH.K_>bL]NbIf2WAX
dL#FKS3Gg:\c8c_<PAIgg/K#X5dU4:91WV(5C\5(\]7+3#C4SR,[PPe6>g:ed@Rd
?D(2R_fOUG6?+/.CWX-;Z4dHT46gKg_HD-84@@<.J@1Q44NJc@EW-4U(@PfYADGK
#CL?6\[8V0bZRL#f_TBDYQ<eTL\DB?aW4aZ(.O,##C=GI5T@)1GG.XEI:6[I@OZQ
=D@Zf=?<Me)<eJSKa=,)>XWKWN#EW@4P+-Y^(=ZMb7P-&Wd>87SZ8R-eg9B\LCSd
8ZX_4X>4\/TJ7BM^@958TUe1>?AK[,;8[CT23:\4YY-?6/CSM2RF#X:B8d54:)LO
@Y4F9EM56UQP>:bSJ(K7O93LXaeK=g;@W3A@(0ef\0_B0-BM]-aB;G/T6_S[GdKc
M6=gd+_]87;\5e6>FY(&,7e\IPLR0<QYabZVO&:09a2Jd9+,QQGc5+A#(I>UKEYD
,(251^Q]A2I\KAJM0R>3EAQeac]O3cXZC9;.=-<T5)e=#_[RB\_gefACF0<D5Z^>
_13N_b[H:5:<CVZ8P]I;YYJQ.(Yagb3-Wd4IMe[G.c@98Xce4;,HTN,75^Fg.Zc4
N/J9E)(F+Tcd/(__gD9b]O4Lg;T3O(6PLTPV)G(?C0K/^]K#WYV;P5#MQ-]TBYLZ
]E43Q1_V2I01TOUWQTX8A+V><D:N4,gS]KHcgK>Z@G;VCY.EV@f.86GB@E/]MHfQ
c]R=U4Gd03@?a#<XOUA<#,U,61@FD1MYbc/bf?28dS>0M)+]MI/&M9AQ@Jd],9Lg
@MH&f<C3DJ[JffO^6:ML.JUX[0b)@UBd84...S5#&I2^c.>fV=gTQ:fcUVVFONB[
46UfG]_;#BRP6g38cJ7F]1X_LL?ZaQcEHX20HFYV^-ZQ?[gTXZbaQS9dV7F;ZN/)
+:gO?).:9=SJg>.f4?eR@/]MP\M5#VaM,g9FT@)/39bc5#49D#&SR[56ZcN.)X)a
YddPRVUISaH<N>4ZFX\M,RS<>>&a=._OJH+CCWQ&8g7.J<_GFbDGT-Z.>PP5J@>.
g?>75V\e<9_f1&Z5O/,+<Yc,O3)9OZZEQeaZZ;(6KAT=M;gW1e_?\=)6\@FSJ)^@
2;4T]7MV8T+QA)0SM(\Y5L3+&-,LH5P[0?7Q>PJ=_1^[K.3E3)8V@8^.YGcXf0a,
&NeDS6;^D4A.)>+WZP3UbGTf+\3[X[3V]>_(FUA5e?Q3&9d&TLH=D_O9a?INS,U>
WHZ5E-],]c@Ec6&HSfFG_I>[c-HL@GB-V8-&VT,Id^IBKD43E&6;)6dT]<GSdE41
gQSASC^CCA0ZRC-99-c(Tdc8#^O?]_F4)M5-fZ0JVJBBIU+-@G^S2FRQ+g2YBb+&
23S>G5gF[1#\I4:cR#88^?-SMbg#9LKC3I^bA#5FW>D5VKYYD36O[[S@P)+a4]LT
#D1T66O)B_N0=,/\@/&QE/UMc<WYNY>,>R_XP,X1d5=e^&.bKC&:U=RS;(X.UL;a
#f^A1=>9^6<dV?b5[GZJ0PR9,8?dbcT<eVd??(<LQ.gUaXRfLYf@L^XYKOL63:[2
RJSa10:F<JAC-gG]H=KFTa5;7_U8WF,AW6BRL]SH4RfJ>eg.QN1^:+NWe>Q]HgQI
(N#/1NZebDg]Tgc5f15^@DUG+W2P\@g@[.Y;+.dFK70+5e-B.GGM>d?1;WXHFLH0
F)(SS#F,UgMOP4g>AdI7T,]6(@3DSK3+YGeAUL_N,0XL+(LDIJ8-<__W]F5geace
f#R=gd8P:J124bWQD<B][C]L=2D9P>a;:HW_+T5]OF)[.8KGCe#JcSX68<)EN<,c
2K[@E7a]K-&@>AD8BA]ER7Jd65XFP=<4?IN(g3IbIDB51eBU-\+1>)cASWDe6?B&
3dB[36POaH,AL^]AN_g3g]XMVW27(Y?U<HW?E[e1#21/(Mc8\_CBVOS>3U.]:b-4
2IHdAP)]2]+:(VRANT&^HZ<a^@e<=PSDPGZNI/6+eI0H(FVf^+f\@F&1\efF:cJO
bC+A(VK#87QLCc&CC[)V)1A&a]Rf@g[YM0?gJ;DM<e2g2.2UVL-.OCYH\[IJe+(:
OHQDL_CCPfA;FeO7B<DA:]=?Z0_8JZXc\:TGPaG-?43NfgG@],U8EQ1#1[D<?(SR
7:XJZOFU.Z34>)2TQ-g7EK3S_>9:_Z?&9ZfK33B8Q80P]&D(a^ML#-;Z0(U-8\6\
GI=EfCQA?<)J_Z^JFg[27_QF=K(L>QV5eb-UeXXX5_=J-_9_g4f?&]80[^G405OL
K@gU&AR[c>Y+DXW[4AOYg7XTd]ZO#@^2?7CO4R.A6CBOXST>HWNL1dM&,IYJN4O_
@[4SZVNb1H@66#0UM\VC[2EHA0F8XXA-]R/=J]NN^fLbG>J_=QW8K3TbBXSOC4U1
V<XaK7e5,,V^ENUB(IGSc/\-NV)>0+FD?FX]9W;,NCbJEM6GcOKV;AT095+0WA1d
9];L>)N2g.fV1=eB;1Ea_e<-(-GM.#JfeIH_T<[1PK>e&D[MYFbFD)060;36^RX1
O_fE.QH?^IQJaJ>#AS.7/b<-4$
`endprotected
