
// // `include "../00_TESTBED/pseudo_DRAM.sv"
// `include "Usertype.sv"

// program automatic PATTERN(input clk, INF.PATTERN inf);
// import usertype::*;
// //================================================================
// // parameters & integer
// //================================================================
// parameter DRAM_p_r = "../00_TESTBED/DRAM/dram.dat";
// parameter MAX_CYCLE=1000;

// //================================================================
// // wire & registers 
// //================================================================
// logic [7:0] golden_DRAM [((65536+8*256)-1):(65536+0)];  

// endprogram

// `include "../00_TESTBED/pseudo_DRAM.sv"
`include "Usertype.sv"

`define TOTAL_PATNUM  1000
`define SEEDS 820
`define cycle_time 5.6

program automatic PATTERN(input clk, INF.PATTERN inf);

`protected
BG6QF\3O<H=I^8SJ_57UH<#-4&_ea9GeKWUc(@PM]b#B>X\19[ZM-)Q-(:^;=f22
B&e_Q7Qc)FO=A3YU.Z]1XI5(OI>[eFDO=#b=O)YNOHFCRG@2PWRNJP0[TQ=/cZC]
/9:AUA4>Db965E-cLE11\[)d_4#U5YQ&U&+],Q-;T+f&H?A3KTO[)X..S0ANBbWV
fJN.]:Q4=I5,D7Gfd9QdCAG^?-FT3Jg_8\M=1/b9=KY?Ma0AO3BZ.3N&VK4#OcOb
:6+Sf/OBA:6Bg_23O7VV0HTc5_-cSIC(]FLU[e8B/T0bgU(@XW3GeR/PfUaW)(IT
(DWd\5V?/ZS\C(:TXH0<H=?.?+\O;QPB,Xf(T)OAd>W6Q7BJTFZO40FX26\M^&Gb
(gM48D(W(cLUF<fT7(K,e3[+b)8OXVL(<33?CIfN3g5_KcP34;H?fGK4NG/DG0(J
M)M6]dMa1(;bF0Ga3R][.R\K\=XG(W=Y3F=\Y:IQD3/Tg.DT3HLa]LMGIF@5G_5O
)K;;;O^=:>]<]L=@A??7XM2:d1^\P?;0b&;bOV?&#N.gY#C.F9^b:#DV0EFSR766
X=3&?>BH6\T,OBXF<KBGI9MH7(N=K<]&+NC.7M:+>df_O\[V4+]:TY0ERYF#1=3H
77[NaYT3MS^,KN2NA7ZBMaH<7(<UfTdT?Je]=LV](EF9NV>4(\@&LAQSc89FZ/R.
GEd:-V2W)>ZT69\+=^-:N6_\Sf>6?,:-<<\U(ge5eRO^=::MF[ceL7_K2D0-)FB;
>R(13=UOaG4L)GR0Fc53(]R#^I]F36d;RN]Ue&X53F=L+ff<7@f+UK-EO:2/Xb#^
aIc;4C<AW0Gg4b<(=NL4M5-eZ)cFNaI9[=9g=>6>?BW@/&:=B9B\4.,LEB=eEDd^
+/Db3-g5T1.HULRH4R<S/88=g#:)W4c[M\N\_FF8c9-Cda>Ka[8\Y1^1-,8ULdP=
;PR6-B\f6T/\M[0W?#NVUQ=??f1(GP<=@L-M^fX(BAa2V>VCKLGYM=Y++5L[SO&P
J^GM2BNN0MH?3I\RV48&6@;@#,a5>da1=OFUT#ONW;UDdOL(6\e3->\Kf6S7T5&W
:gPD?:D)2YN=egJ\]FAaGI88gY?K<Wc#]4@+C[5.QYHVRS@\LM.6P)A>IB[2KQ8Z
[_0FMbdAWXAg=J8DX]a>ZRd:0J=1VBP-7:](]2V7FLG2gQe7)/:_6R9(@50<]5^2
[@GJGZX7WE#[I3Y<aAc-IU4U1G/@.\THPeX:26If;=<78Q9YRFDG.Nfg5XQ;3B6E
3d:f7Y23#=g:RKZJDG;a_0-I3gIE?2[H2>#ePPZ+-YbX^;+/9O82EV/a\Y)3-ZL[
c3&d,8X^\@^PMAEVF5^8Cb],3)Y8>Lb?HB(V62bU9CEIGYDQ1e[O(C#Dg-X+T)g.
ML5AWK/<CFa,G_)JfTJM=AFA(P#+]Lc1Be6E1fWOWV9>B[+#5=I1g:Zg2W2D6<N1
g<F2XdYN159dLNEGc:C9Qca9C;M^NMaT>6gYL4_TH+ZZ\_PeO3aWc]eKPA=1CO\1
RBMI]>AQ)X491cC9,Ae)W8X?&f6W-?(U+[XX7AN81WUZ\Uf]&D7VG4Ag:+,PN[:S
PLcU5#?CGYJU_;OJU^@507):<X:(JfL@[P5EWB(O&Y4)^b61^cU&eU@SOQ5>fS=X
^J-?Na,Z[I#;6JFIO3@g>#7ZQU:WE0BIZ=4e?JVTPG/<#(XO:&:cA/#[(3^UQ+,W
]LMD7T@cA-D@7Qc5\Hd?4cGY)B37gYa2Q4^TSU8SJcT#9Y]QA.d5fSOYaeNV;Ig8
NU>CPIXW7\6@Hgc:+@I92-R2M+M_(9_<dW4CMDgESfO^.-Dg2]<BU72?A_)HV(OX
5cN+34Md(L:;HJP>)b#L0=/Uc&fYNRHUBT)=/UYWb/aB0X\?a^<>:?SZ?6RIeBVX
69\1WFA2QJ4E+cV[=S^QdQ_>\IID.c_+3,;+9dMSI\AK.[9d?FT_8X^2gg9MLZ&>
VGgCN8_P^R^3M2?U[QY7(_TM0g@B\DW7b>fB8\#Yg.5=AD8(QMX]/Ha5CO(1./-V
If@1Vf_<,NU^QOPLPb=7Q0?&6Uf?M\a9-0\JdeJA>XWUM[;2Lf49?HG8,]fWHUXL
#>&T9a#S+32]8))J+5KBT/-Q>Jb+H^+O2M(]d,N\J1W^L^L&9::3>FEUATfGRI<X
]S-R,];_cA3=,@[5OXQ4d:I)M&4S<OVf8\#;S2S#dY.cE154EU^gFTd?<;0QDQa^
4]QOQFF+/23&fOI]34XN(VO>8SP0A#QB6(L:>Z,c1SX/23[fEQ(KSSL(fE.5;D&/
We+FXCAI@-H&G8(5ET:23/M3ZW@I.?^U-USU3?#G=-TOQZ4Ya))NUQR?Yg2C=[UK
JV98.:ITHg&H,:/#=3dPcRKP(K.N-/4L8Xe_;D3?@a(W30IZ>=cHEH0-TEI]WT4P
RD,:[[-A>dd<5)FC6[F(BZ=6F:?O:216Dg+U6dA4d(3ET1,e&,?.Q3LH\RPZ9A#?
Y]N_DZ-e].PIJ4QR?77-7-X[W6XY7g;f(Z-UAA,IJ9Q2V+BOf7K7bVb.f:L7^0g)
;3M\ATT#=6dZFK90bDOL]=DgJCI(L<SV<a+A>QbOL0U:HBE..+5M.B8AU\b2.gVX
>INVO1YKEf[g34^KGUYcS;W++S96.2Ba1TETf6d,<HG+R2&e1J5WcKN#(YaL7_3]
KQ;XDgO\dODX;+Gc3VReb,WY,FG,Y&d)9#WXWQ&&M4CJeYS+4eeEP=b?+#6bNSKc
H>a)/]QXP03KU([HAf+^P0_89S)-Yg5RWOgQ)W3M.81F;;JV\=QD_@Z8ZB+9]ZS&
EXWD\7f53]\8#[RE-M/25\RbVJ4\-dc:]@YPOS(>:TZ8L)=F-EP3QL2a(O#FDCF<
=ET0W6]KfR#,@Vb2G<6&bK,/?@ddQ(XST8BD,b/1=CY6ee9bL^7,Ug1UcT?;JE[<
;P5]YES:<VD:a@_6U&).HS<&PHOQAbB)42M4>fC@5-fGbN?VNB((]WgDX_N1[KM1
VGM9g-6?:gKI=]QOa)X]2Q9<]4&eb68>^&HLeWL?.KA4/5K?]6:H[5B7B@a^S9YB
GY#/C8GODE>dX2].Y8K[eUSBNe5Z>M^e\XXXRUQ-INL9d6S#ACA.(K7H[;17F,QW
9Lg8I.X+b-R6#Qa1(S1aK]dP9e41d^/+I^I7FX0BEJa]-Q(;MCSPQb7<[B2eC8U-
J\6>J<fHC=XD5R2)^_L/NL[c(DO4BC-9L-XReH4bYQ=9\P9/;B=eO/<f[bP<=MWL
VgQY(]9^JL;J[NYZ#/.AS52Xe,0fbfJC,EGY^g&6bIAd#Pf-MfK^F>0e4S/.<I^G
f18KR=:O.IARd;KXdJaOU)N&X<(MH.dDX#[XB\X#JLUL;)c08#a@HM^]^#U9,(+:
Q>B)86^C\AUZHY,^e2>,(c-5635d<QKN8\8_N7_-VP8gKE[cN;f@]YL;bP+0_JMA
@>dG(/V3FU)C3BJ_I-]R61>#F@>f1@P<@<PB+Pec2CO[O()b)SNcAfZ:7Sg:6SR1
W9:<eNUdgA.b8YSEP6N<Z7?:3#eg&X(J7.S7-1gFU>I<P2C_2+_HEL\gXYR)bR-A
_4VOQ-@T@cGK8LY)+Y2/7gO#2<7(GO83?&2=6fXdL4+SWAc)2^17<XTU[GT7N<O:
+eBHfbE?L4=^Q^HT,Z->ccSR2LbZ@K4.&:4;QGc2/Q8<1R3Tf1[)0&C=O6SZ).bE
L]Pa31EdOgK3gH)Q]RLYKS;A2PCMMCY7_-Tad(J[.g;cLVX1#U<UJ=Q-VDKUTf+f
EX3N=ED]H)aJaPS4;-;gB(Y</W.Tc59IZC:;9?^CXc+9E7/+VVMg#.2.M85V2DR6
F&7YJ6eF-c_Rg:cQ08E<S)OBI7,fM^ce.=DS_8Ce\WFMZ[2bR6VT9]\Gb#5JU4JK
TO5MQAZOOU<3S^_108:c;2b7_AcWX\6/2C9GIF5>-W(,<6X26,(GbM5?aeQ.M_10
dEB59>3fFB5c)TT)G=@S=]eC3#bU2C_RT1:P#7SCHL9@2HPQ2H&b7aE4<47CIaH-
N:H(L/A07F@Kc7dIb##3Q6PVbPa3C#OY[G3A(<e8ceFZgUS::93ePS]I.R@IJV11
)_./L-R?6CAV=OP+:TQZXe6G=;c(@9U+G(8=OR?_#P33]A.FgaYZ(F2B0>(LU8&J
4Q2GB.W&2_7RI\]Q>A0E\QXKUe44LH^&BaO8EKH.:8f/:FO=bWXXF=E+6YNJ@@DO
C9H8LN_#/KWIV>IcaKX3gBc0&I#&DZ32#,)2V,J?LcacZU-KU:Y@cG-G=S(b0+XH
NQFa7eQQ#EeJC98f>12aJT8)Jg1E&(eXE8VbBCPXfVd4\N]G0fc11dUd3H,GR3CQ
c](Ff/dI0bJ82N;&6299QZENE)DEEE_+aP;+Re/c6M>H\PP//8N\7cWF3#L\0+-P
Td;^FRH7GJT\W/I7?2@9L7.RR7Qd4\54@B;L7WL?34bHdGMcX1Oc+g)57QdW]gO1
&b0&9aQ42:(IH9Id\XH@(]9FS/Ia7ULLCWZRNe9g]:6:aL=X/Rg(f71+:W.PD.34
XWZ@=Pd@M:-[8&C,K^LBR_JRFf2SU^Sd/f.-P;H@N9e=BMg+7)4I<]ZEaUg7CeET
f4;Z9g6\^E6#=F,VaScFJ0W3V;_3ZJ(F-RN>Xg7Y]\_)WLS:aHgdWDRfZaJf?/f9
V:4M(SP50.@1M);g1#]c\EG.gF]U9=7ADG,UZ46R11f9E,7;5;UC]WE?MH=6R1GR
JDc^&)W5RfB5=EW<WCJ43W<eTPa^E#B1RH4D^cP?21#7SA]]OB@5d2N:TGUJPZ_E
@MB<\L7>]+Q&:<gJ6<>9bA+LaZJR+O4a24\8\OT<TY[)O[+<VT<)[M)L9JAUc;IA
5\[F(^LK_3DK7>=d_e256Z=U<1K3^0V+P@cDg+Z)#O_1-^G&?92)g2XSGc8=T0[3
4R#VAT)Bc01SZF.T3]/<XNA5S>,22U@f7U8AP>]2P+CD24EU;R^:F[#),dX-&<T2
VD\ZCXcQ2_YJGO5Y)Z<B8IW9CL9>@1,&;)C1;L:>c=PFeTY]F9GU7Y/(0M:8E5==
I7Da)VA)Z9e4.6\F(R51/Bf2M]/aQ47E7V3.VfSCFM3KU(/V+_>+AK)4&&JCQ4X;
647.B^LfX+beIP>ZgX/ZY#5EHI@G2_8L[VFSR>N]C57,-E^UL<@Q;TfJ^^3BLBGL
<&\-/#YO^g;&U#<COYX>]H2^UQbV1ebOR[D[.#D]V&CeHD?b.].KH?e/<S\V-WKQ
C2Ib;XLT?1D9OFE>N;W]PREQD142QSR[M0F_AG2DGH)I;QZXJ/_[D5OaRFRA1=]K
ddaFaQL>,;C?TZ;6U@RLCe][aU&>>&A#9W2].,MD(JX(0&10<PL1/OJ_G=_Yb0Qa
(D6[-+?RAE3effU02O<MP.+9H5G]6Og9Z^DNR9.@aHK0cKZbN&L-_[JD#-LD2GX_
9EAIO^R9&f[9>HdW1T)0@=@T.G_FeIbE)gQ\P@JMKSA:Y9&?890<,O6,0dJ0)QcO
(SE7#c(>WXN]b?2^)43K\>M;@J3>ZRA9C0HTbgPHe56^d\<NN:HL6Fb<b93U+@YT
bfSIa\[;YdW/K8E28X2Ic(.=c4WTN_@KVH/Q#O5#2K4e+@eOK);B4S=3#P30(<8)
Wd?5+\JF&Ue\JW/N=3GZ3E=7>cb+ROM\FA#W4E>eAZUG^#=?8U)#bR>[R]CEU5B7
6Hd13Q3H3YOFO&463YKE101U_@5>X&&^f??&VV^^#Ue[a?R\[L[/7#ZCTEX#(I4T
CHd?=W]J)->-Z.]F-@(N]/=Wa2V6M:&\.Z:;5AZRI>&OOO>>Y84D,M\_[Z/9eV4L
)DX448S+H;_>Qfe6/f1(\);c<&T;4O+9Z64YeO,^-N>]#9.HfRgR>05=R]@@.-JG
ZDNK=T18GODPa##K28\[0[RDHa<\D3]TE2+c:cAeVI=\>TQ/6X1eZOU[#/@cE;MM
3_CAK@2N2IKE(8;S&eS4g<H7dGX1,9;0f.EG70(SVa3baIER8acK,^5[=b&I;2YU
O=U:M0#JP)3D13H97ZU^L).+N>-U\KO3QB#>]Z3FEWI/N[D.]g3?[-6LYS-9(EET
4:fTfKF2_[6]C[)?d]6V.^MT@<A5;.a(KVD]+Kg0T#=aaF5-.+-_-Q_.L_T2[W:=
,U,V_-4+<@LTF5<\Q71UQc^9V&gOWY5->^.<#7fQ@CG]G;YWE+PD-[);^PH@ge5g
T&U-LGMMF?,WOMVb06+&O+#SVU\+3e9O<FLRV4XB@fAeU@QL3,7J+@@RX&N[F6eN
gV3I2@T53HF0.CX>=ga3BC>H=f\4W0YE]b2E;6(/K8NUG-]93YFe(,Y>T\BdJ?Za
#-6?&fEB]bMeC-/cCJ#dL/=Gc)SH:/A2\3QIec#@_ga]fN?F#1719<^2[-OB98YL
Cb>#+>/Z&6.8?A6ZR\Lg\cfZ=,NY1ONda9:8+7dT)f2QWRg<]]&&TLUV@9][^Leb
/\NQ2/R8YK[A)R.8c-31@_@S:f7J4L02?0CSERSU_dH9@[+,388Mc.HXOJZ+57+)
gROabSbAYU;3Wf92#:bI]+WTPU&GWCY4Q)OOMDCGL5:AI<PdNR&E3590;Z2?I0GX
)_6^>F:-VM,6-YFW-#J:5:P@SN:QeQCR-CM+)D7>QT;7V37HWRZ;+TG/SFALfa[e
MG?J+Oab/Q>&.91bR.-=9;fceOa.=]U3?VggDHI+c44R].(PIbI<BS()M(Eg>6QM
c5SK2c9^<9G:2LOcUH4JVe9b]#?5PN(#<9>3dBE>52LFCWV3B)Q&fCR^PALV0D[F
ZZcTAM+<.BbI7K4L7V++:YGQ8b@8E2MEZ1#g]3d2QLX3](#_e3R4X8)XaD0;SYM^
Z?&IP1aNd.4b;Y(0+T29.NO0)<S:6#fZQ6f3LMV)7#;g>J]14WG:T^;N.0Z5/73B
PH7</_[B;W\Z5.^L@CaIa2[S<STcCAVKAD7</N7;b1V1SAIIL^P(0aI^<.eF]UJ8
(<fFK/2<1#W=@=AOOce6@?M:C(<)^CN1@@aa4Y)5?\,)P@JB6A;+6add2RIAgc\T
F4OGAUf?;:FS1U125&LUYDLMKF33G-O7-YV?aA[eL##K)DG8)6S2_Y/LC>ON?aJH
H(:d&g1ad5aUHgL+@N>F^X([e(Zd9&&^b&e(/IXYVV<VX8_@]-XJaR[OT8gOWIAE
SGFg]f1HY\3[.MZYPHCg&6Zc7M#ZWP\]GPO<<QMdL(]&Kb3b&0WFSdLOI#0J7IGQ
I0A]MV=gF^A0WdS]QPYFcGJCZJIV7SU5eK+?Y4IW?Q\c<0&EZbM1Nd7E/d+ON79R
CW(2,cVZf4?1G[8>b;eK20KbS3=QD,-VIc/YW?Z@0430^V@^UQ2QX&YRU<G)?LKG
Y)X<WH6Q@E_I\^LJ[:1@2=.\5g)<4@ADM+1)F)Z7D#6.8M5E#GVgf1Q03F+Cc\[D
/b3\Uf.:\b4N:#d3J9ZJX6dF,J#e(c.C;,;G6VBHJB8c#\gKB?4=J8CSNGERD0Fd
c6)I_A\9LbOf4cQ5#RfUg&K:Rb?3S(T[c]_A#+\Xeg5Q6I/ZC=gP091g5<JgQ#/^
GRA9d>M<^<gY]f/+,=HFf13+4;Ha\0Dc#RgT6f4>a]aa_=b@P@(W=5#]B]dD?a&S
ME-1M;23N,Z@H<.E+2d>TY;Q7bR\&7gecaZUE+;Na701H/B5.FdAGc0V?.2]#CC.
EG6RG]C8H).UVeD=#VKUAVM5&RY06[ASMKB:f&@ZdcgIBC[:2J\ZO:.NLWX2ZS38
@A0cb,VKdBaOPdcP[2_(?/H)V,[YDV_d[;Ad&_@GV(#gP.D#5=D,^(D<7eP[@<7K
C/=g_-BJ-PQ_Q]bY9W)52Y_D4&&a)>?BJ.HUCU(P7CIW,QM2TBG^/^];LT8_L[cB
Sb_UW_+D>XU.P(d44GT24D_U]EP6UL^](A6;QW1VIWO(M3@BZY71aGfFd(XZfQ2V
]O]c&/49YA,1YbFF[S7TIF:AT]L.?PVI?ERNGa,P#@^\LCW.Z8TUMYXa0J[2)3JZ
:^TM)V2Eb+_NY27/_QMTb2C4ZFEdbAACRWW3#:W)QYDM>#W@U2QN/=gC#_F)a0U5
W.<P.XG&3_>NA.2c)A_N4.)dQDZ7D?1E3:U.+;eOGP03eIUP,.\Jc1D#\P5d=Ta]
]24/V023O&O;M4-dJf6>&UY=:M4d_EcE-TTU7d0[>=&EAM899X+@BY#;Q,^KC3)9
D7BOOIfR)BH0_?eQF)PY0fgKBUP>YQH[\-,a6T8NIZ+0Q8.1Rc_<dZ>ZP8X1F5ZL
SS:HVFf4>4ZTg#9[M^WfP^FR@=>&4QJUHE&N3139g2;?-dSNPOFA8KQX+37AJZS^
[LT#3E:CfV8E:TUO.-;NRVLGg3Y-7#TK&aJH6aa)TG3K5ZDMD3c2I4\QA#T#gO2b
=O/RgF05AJII;#U,>b.NO]&.0#V^XKdc@[.?VA^f=QV6,S[D.DBZO-D,M+H5f?Wg
G@QXcE-@,76/L/L2[K\KLX-H1e)_L+GNYT_BB<7LEZg>B0]+0&E&)FdP&YMeX@ZS
<LKb1Eb3T1_;Q6bKeXV0Hf]57;3-7[(1]<X[9cCd&8c1A8CZc)>O3ZMPL]3P3ZZJ
MOdU.M>e^8YbeIdW-\7&U(I=GW3:NGA>\Cc?#EB@5]+7BE+@@=YF25L7\HWE-5&\
P9(8ZD^/P#6Hg<Q7/#L8<<40I4fI>ba#fGBVUfT@4b/d@U\3)J,(dS3H+?D@:#ZY
dWV=V4a57K1EP5)^[V<5Q_UJ=>:/aSC/YYQe^deYTFa<,(R>1E3>1DY@A//<a@FR
6TB@EB>0cX1>d3(]&\MO3Hc>ZPg3]dQC#b#TZA:V@f-2g\K3dFNNF6JBUCB);R-X
DM+<-/QMRL_@eGd_JK+(GeObCDUCf)f-T(,6D>W#>,73;;c\?J8Ue(??d^c\&dHF
&PDf(&6XG#-,)[Q+@cc5Z>Ud3d,Q:A8:9FA,/H@/PE+UBS;I4e__8c\RL5F2EIQM
abY>YUEWVZ]BH,7J)5b>g391VbG0.DX.^H)6OZW9D]Q>WA0Cgf^fHfKRTg[A22X)
c/GD&VN<#(YV?BbP/ZRB^I01NJT<9-]f9AFdSbSeGaY<RP\I<BMDUHRL5Bd)Wd45
;;4g)RB8UBPN&?I(D7KI>c?4.^9+HG=A&#bc:X9SSCT1EJfeg^ff:E\QKW@<0OH+
[4&<8Cc_T@WZBWEdPOM]JKS(Gg\ZU25A);<EE73b,>,CHe9[95VC[3NGN@JW-LH2
0EdZ^H686.5=#+]@SaCTMUIENNS.g995JaI?D0]#NU2Z8,@;C]0bT)^5V/VX)FB=
VBY?cJ#ZVW;G^;:7WP17S,LN--)MO<,JeL.]:_;W_><[7g:eYg[5..G<HD5Bc&Ue
AK_;2K:LVMRW>B/5B]Q4bUA/XMD-C-/dPdD(gC^<^d81G1[OVDF3>6B3EU&MJ=4^
LR/PK7T1=aKRTa].<MHAPRW15]W5(8X+;DSS>ecbT30_H@<M:?#e+N\fK91Q2)FT
TeNQRV4Bg6E,8\fc50M#^fEKO(;?<N+bVe&:DG@&W;<6:GN.QN[c9]a@,,<XTZRN
7B\6IU,428a1;KCZ[:6b,3N7TQ7Sf-A7\)D+I>Q;M^cVHKS(_(fJJb#7N2H?gc>>
4?P;G]X-1Y3WF^7afFKMYeQ_+&aHS,eXXE]0gN:_WY8JTbbgDAVgG9Q:9.C07<G@
)SCDa,Dc@F9ND[LW/Y)(V<RgD^2eP8W=XL<d,/2:fV8<@,>4e>^G<c7@3/S.W\D5
7ENK&44)6ZTc)R6?5OH<]2_OJ8F2;FU0YF@^00,;7ZT)5/Qd>g.7GM,5gI;7VDfJ
5@_,d?EX88B4g;G?>?2ICP7We:A-BWUMKNb@_-6e&TQ<Oe<#PdG^LNQ[WF?8EGA#
6(HEP?LV<G>J.-A.4I9gFD:?8cQDR=&U]&N.R5Y(L&(WdHcHV7/PW:]a_#QeL015
JWS1\T^]U-Pa;]3/25&AdQa/ZBE4LT.JG-G2-c2NbgQHI>@W[_cW_A[+5F@,;dOR
:J&TJRE9DAFR8920b;W?I17N+<gRReIKA(IOXfcX<?E2CH[fW\Q<V:7HSX9N&UGc
J[>6TcM:A?,>:XRHc?LH@73,OSVM#:SLE\7=4RLTe?YR^4A(9:186VODUR,TZ#WU
]3V@ABUKdH:gT&>]gMW#AC_aCRRc&XLJd7KNfa8MJR@FD&Q1a9&<#4e-[+e6\KeX
RD_[#>WgPaG4K=YI^(+1b\(\L+OH^#M.=XDS0UgLeg8(UU2J>#URPg1S]#/e41VQ
.\,+4(4T105U3a+MMbA_SKCc1=(/e_-510_LO(d-E.@OE.SH-#GO)E#eVUJ5aXA]
CYYOMK@_0YGACRPJDAcMB0<HZ9UV]6(+25Z/P+A&9<()1+7.D;de7Z1MU_b#<aG\
@DAYV>J2[..)=#,T[TA7?_dAA-QY(J41ae[Dd]Le<QO&;30=BI@[?+c(R2?[516Y
7D1A,5U0KK&b&@@,WE(VBR:MHL&AY.),@,EO5BH3SWcF92cLcCTU=,@7)[JV;/M]
<Zf1BFBHRM2/a4=PJKEQg,2422(<]R4UD?-JAE)Y.YQA.eK.L80bge<;f/a5XV_(
34S)eb=WgAWZB:5<N+YHKPf/gfWfcLX>cce]e3_AIO2&DbER/E/K9NBd^LDa3TQS
5f0#XF-e9,dLD\9e83/eW]--H=CJ[X;89Qc0IHFGcSX3:R_EPgCA1d3[VX6/7I11
7ZM)f@&M1CgW0>Y@P8)g^ecOIPG<@N5<a4X[O<P93G>.1Md:+e=,A&YUP_RCE8T4
<d3;e@PCT<6S1SB9D#T>G@M1dB_2@,[>@(dW&fBI938&[;B<Ge@W+WIEef(04RR2
FKG>008\?9=PcPY9+-0&Z-V8,a>X6B)]6IH7>V.&J;9E2d\R(XP)@7^<&3(0FEDZ
c)Yg9+(/Sf-/^=B\J=LFF,<6GMY8W)e=54e\V,-L1eQe&O30_IJ@D4VYWHbHWZZ#
WfOM+ZBI4XZb(Z2EbR97T5d->^,=C<\gX:-T&CF-;2TA;)RV]BN<S:VI8UO5&f&d
,EeWES]FGa:32=#<.;85(b[7b<a;b;;SCG1M.Y(c__8I/XB6ZP?\X_4Q2PEZ7/Z1
\2_)35.MdL@McZ]JHD6^+Q9B,#G7NeIV@1eJHNAPdd54Y0HHZK^;9D888GX=R/A4
1WaJKUH,@fVbb.J\[L[gX.)RaCKRJ5,9,S^=;LZU)RV_a]J^<\&4\:gEJ4c&-#[4
OHL<@@<NGEP=TG1ZSX[I;@=EOW427Q[;,@E@6RS<LDbbRb.^/5&I+03T1V,>[6FC
_]K.[N0VK10<WOGV5I:gFZa:+SHG^ID:28&G/ecN4<U6J,6G82+2MQF&@TS[TP3]
+,_Ab8&?/ff^Q1K>EcOVO.QS0QW;PTW.1^;R0LS-FS58S56;2S+79AP#I\)7@4_E
g<I)I)23Mf,caTBc(X5FHPVT-1A=11(/6d=.c_P)M@Q/0B0bXYWg4SL9=2E2,(Wc
\@&JS)&Xg9QDB54_A8Jc9(;[50NIRQMVIN)UCV#]Sb?>9>G.aIK(=#,BU=IQ00dP
F<&7#L-==Q.<N]eT,XZ&=6J7DL(C0#LSJ2W(;GTRfa2964cIgX1W=49]a+gFT5K8
Z,93>WX>Te;(1[gYc+.Wc0f78QTb3-2ZcEH/:J=&A(7=4X)\G^bU.,-ZOVYI6_\L
e7,GY-GD88J5K<F;B>(ZHPSTQ4VP\cEKfW?X4^N3?4+FI_Dc?dO?KUV:KdT[2[TH
9&7ON#;ZNfJF4F]Y&X,e[b6+7aM/WXLOZOQZ85H32IQD^3#:#c1[d79CbYVAR/X)
ZbA:)I9[RQJO6YP+)P6LUGQEBZAV[20_L.eZX_B<,GN]UcOCN\Vf42]/ag.4Z6WK
f+SHGVCM[Q>+VfE9SF]g<CU/\YJP,R])H?.H3+<69032ReQZ;UG\N+11fTdB>H\+
b7b=\@@36UUFQDET7^O5PBC?#\:E0/=V&fA))5Z[dZ9VXBaQ7TSeE?UD)@S^#+NO
:\7E&d9;;0UCK-7fHUMVS5b;TG=4d#W>9<9@fD71I\4;TG&e5H3d,(aU>[AJO6KY
J_I/R7:bR3VMDHBAREPc=IDBA0X5\##=#I.)<Q#/YEIgE\ZcH2d77fJ-;RXB82=+
J89?65E9F(IS2KVM].HT27II&9&M&/2;;a<2@gbed_7510/8]@_Q5C<=\O3D/A12
@S._@3+V:M\,1P)A2<X@\27VR5MS>0=9]Vd\ceKL>0#J0SCS2E2c/RO:b?[ZD,Z<
e84c(U1QfCPHB#=>\eVEO7<daFV\J76GE9>BM@2e;UaCO+5&Ke3dZVC]DdbK800\
0=X7J;V<.8KUUV]^D@1d[U#\dDN#/^/&XcT9R^^Q(#)TYLYQJ63U\&eL@W3;Df>U
50M[7(_IcVMJDB(c]KC;58gVXQ2Z-[)^T:EWF7(bK-Z82//EIB2FMfPXU</6c5V+
dAMRZ<Pcc+9-))YO60>;Z6UPV2PRSfFW@_2]69Kf,a.L._HJ>cc;aZZ?[G-MVPa+
6KBI^/YA6B5KL6DD-OdR9Ce(.B>-88e1A[AHW)\1HJW-0B&f@\-KMY[d;5_5GcfD
6=@+TROKG,LO&bM[24D=._a.;DA9I1d.5fdG2WEF,]4.bc5>YFN^]MH:(f?0ED)F
&eZ&>QB:P&PcYdb9ONW8Sa:,:..EO4JUKW6KMA=f+cL;&)<MDF@RFYV?BO?(N0Z2
bD5b^:0\Ec_2HfRFC<N8R5H(O^C\gDH2>CI\9VQaZ:2.aC53+P5/UC#WZ/1TKgN<
M/TLF=OGQc0G7ac<We4>JEfd5gd,F0?gJeVZ43,a,VfFD\.^=H-5,gSc.4eD0-c@
C77b)FCR\c<DUCS[&J<g+.JE\K48;G[d1^9[1.be2a9,HW1U4KW4SfPAa6-P(d?,
JBW#fd24Qe2RK1_/#?N1,))6>()E730I(-,H8H/ZZ^J-c@?XJ?DdS14X5P(=d9H=
BbG:.ac&8gYI\Y@6D3M@MVO/b_LL#ER9Q32UU[_0+G@\^,RNfA;@S<1:U)H_#K7e
R1\bfU6Z4.)_-g-Z_=#.KQ9^VT+(>241X@GRM2OI9U\]>I,E0XA#Z&IZ7_+aSZcO
KJW,K-Y0f\F\7aW]B=B8^7F^E]/O+VH<5\Z>d9eFW;BNJ_<>&gaC];,<F^L1Ra&+
Red\@RCaT<2X)=TaHF[,e03,UW3R;fJ-@b/<V_PaKeIb;.GEF?XVBgF<b>P=<C#O
()K(P#aP^XQ7McE<V9@cN0RT5CPWD]XJR-.d7Y>09XIfZ<4UDC80H/GG-/1QGK\]
R^GR.H9>^9=C69<[PcV927H#dT@FMBeT34,(VXFN2NZ<<<+YCMR1b0e>A<\I]JK]
>FdeM0N\1_,?e:gTN3g&<gg(2\A&KPNAZ7KER.?C8W4?De.BO(]?BHX7KTEJDQf-
<<MY?-L(^A1HF14Q8U;QXd1EJNNRO;SXST@V@9?AS6Pf/Mc)XZGD&[3#<WZEWF@/
S.CUR?4R\La0T?/C4g(#/NZ_geUagBG-UDSP16WL.5__/e3T]Y4F-d]-G@GLEFKD
PU/QfVOcgNWgK:f@KU?HgN7dXbQXeBaR<55SH]UVKI+>@fR6DY[H:dB]\VX(P-],
V+FHJIf,Hd-OH;bA#@F0@[b5gW8V1&cM:d_5HN(CQ/.YO_dQ.9),GWI5&9aB.\D=
IeYO[+3E4bH^D)-XA^V?+@MHS/93#=.5ObB\+-\0dNOGfLf6C&E1&-WdI3dSLO0D
0]Q#KCZ#<,>acN+>A=bF_;\LY7PacY[bK&:34N^[R6g1_F>JU[Mad<OL4UIRM&HR
Bc-O)VLD[-E]J3FP/X\PgY_F.(2<PPR[aQ)J)?a-821A.2,Qb;&+56>3#<47(2<U
CE_UBOf@=9C]=fR4?AfPc_\JgJJ3fDb#_UH622RJLQ3:1#64MF5&FZFeDWZ1OHf8
Y[V<e-9=AGdb.+A)#a7:>^+1dXR9e[RF<0(E,58J2M[<>;(f23@5E9TF_TRK(;[7
5\E5#a)Q<Pf=H2M.RQC2P&8NNf9G,@;(^9]CFS0-DXfKEU6Z^V<g__)\bN<gEFX;
0\@:JY9AMVMI\5@^?9QgPC7GM<aEQHcYbY.,XHDU76J2L/Ma2g8)b__3EOag3S[_
_D-92&Z@a-7aP9\7a.F/L=L3,-ML?J.WV6bg&gZQC>:f_K?[33I<[96P<b<O?[14
3/KJK6AN:&J-<PDRWAJ6,edW[MH\:28ELSNE>_?GFXU)2J2bDXc\/-V=IAF-.II6
\D44(&,UNK(bd4[N?BVef2]dLR\V_O&dU[.2:GKA&35.)SD0<@A(H+I>UV5>/W@#
F;e)Z8FX2P@OS+9Q;O>Y52\U3&D&[LN0IAdf+OK@-S60IQO-L[_OC[WNQZ(V65JD
=QDC<ebQ[/W9dPgDfE71d517(:e#dS<-KK=09#IISB-G^[(+2fWdU#:dL,E(<-&e
R#f;b-a-=M0VY724OQZ/,4S/M>5V8;OJef0#g,5A+=@D(Yf=_@/TFY[DB^G)A8\,
&W6XbXV#YaT,E37AQV.EdWA4J.U3Z5^:=E3&F4GW\4XaYVPb+=:aeYD((-gO#3Y9
G4?GKGgO?MP_FcTU#SVY]_4PH@KDQT7YONZ6\aQ)2HVK1/?.;RaI_g7cL<dHE<QG
1SZ]gc4B#IALfdBD6<OL(:eROPcJZ5Q_QN/a^YPW]Q?P@.9KT,fG0B23d)2OY<Xc
9V?I?\//4G^=da1/6&VZ4;Nb:&>4(C<@2UK[C;OR52d6D6_8>V(S6QQ25@[8R]c)
;,7>BJ()LM^5E[cK5UTb+;eL=A6@dL+3F9cJOKPS<T7dN7N0G>]MJ@/(;MJ9eTbe
#]@W201f>.4cHBfgPCa,PZ<AR[)KePZ9Z,/aZ]OU6P0EHQ9^/3eUaB5gGVP1VMN/
(B=geY,S1>70B..?RZ9&YY8g=V^g&W[2X5RFX1?f^:2c0e/L<VVJ,@XLM\),I7#c
#g1QS^,FD)V/(Y=,MGf>f_&<KE5dXO,<dJg53J6.OTJ#fMF^VD(I=gAJWP&FL=/2
0\[?g<fD\ORG[R0g3XUO4af5:cd,0Me]]W]E.9MCg0[:^aI:Fc#&Sa..0Xa@D2]H
\5(gCH31PNAg4f.aJ5;YBI8?F>eAB?V.U(>:-8c<PWDN+BML;Z0&,?PWMOBW43IX
N5HP&\.>EQU[J+L/A.LN9C,>TIO)J1N2A(8=N5\d<J+@9?#K;)b?d2/dWX]&cN>1
21>d\2Y<OA#BV_.)fgDI0INb7ecYOLT4)X-@RNILC/B&W,]1#F)^F)0bcA_cZZ4Z
]1JB6SUXN)WU43M,]H;@E1]_NOX]TUd(M<=2ZWfV3B)^fD\)UW2E@HR\&^2P?K7Q
\7G&+ZTS[T.(Kd4[<79[A[B)aZ?FGb.\G@UgTd..36JZ[A/U@&N0_>5E)1XJ0K-3
#L.@V[:;+8<+CHN/caLCGe\ZNCZ916ZV-]<D(_-)<M=])HY_VOEd><4a8M0)dX24
UE+=XX?TJI>H>XI.gRLUcZ@Ia&LZ7@>MYX2>EFTYOGYCM-5E@(e2c/OH^.ECe+KF
4(#I6d=W2O]=@),DLQe.Ea;HdJ8GRYMAKJc#49VNY8,4(JHP4R;?3OCH,IUQKgF&
T\4e9&LcGHMBZg>_RVfNUTf,X0?gK/(gP.?)#,Y(&N16&Za<7LWdeMcUXb;[9RgM
AbJ.9[6@N_]a/RC+5]16YBP99SD0P_EG8&.d^U3P:)IBb\@93\57,JLL>KB/P/fQ
/KIb2,X^g#ffU[#Y(N:=>PAZfH=N)FeWE?.R.Qd?CK.b5L1-VT9cA)N(@R67UI.8
e#Z7I2H)=bd#W9(GYBB6C,.NOB&eQ1RE2R[<Id88UD\0V>@f^KAG:1U_S)X77MdH
RK.<;4G?_I#K8AQ=XMTGdE^V8X+XPE,?O]?GL>>,a_92[ORcQR.BFK>.Ta:/X-]/
\G>B[BU+Wa9]F:XX96P9,M6(@VJC0#V(VG&R[CB-fReA]LLN#,6c+UV\,,[T6)7X
M[CGgfSa6QVEL@J2Q)/K>5]+#@.N/aFCR6CQDfO&9C3KAICaPF0BLK)?=C;V>HSH
@AZMJL),,/H,>,2bOOb&S<aC66L-578;FYFK]F?R4/aAR/X#2C3bHeK[X3SP2^b[
_[PPb>TE51cT:\C;?Rb/3O170a0,CUe6Ye+d:&Mc#b<YK-27#9)N;a5]]<D-87H:
SaEU4M:.K19TCJJ1a;Q_;b+3V1:6bb^dbXLU_Ma^WOFe,Q@0R9fF6aU1O^H.b.28
3<-T-RH8XbA2faJGI)02/3Q922JQA?8;g9)N\AF=1]_KcgDQ:;/Z.GSH@O@Z.1ON
:U5&/+\3:9,I<8+O6]W7[\X.Ee6#E03fEJY^Yc=KWb4I;]d8_K@L2Mf8ROIM2dY7
LIeSL_YO8LAY]LMS##KN(,L@QXC:/B.&:[^g6TfA+T4>V#/K>Ga#b20W,2^eN0cE
/0C=f9DYW,1?0?Va&+)[6GgJ6K6@MfeG.GZOd\-Oa/-gF1aDH:XXG?:W+eIO&(=P
=HFZ5^(TT)4C,FU@K93aU8)61gCACT7,]=3UIQ1aKZ+:QV:b5//@d@UVQPQ\Y7]K
d(74GEQK/RaU48.^W/>:baB^C-]M/6Y-]E6&^I]5,fF(Y0A,eCRF^AP>1:,b\T8K
8LV]BH5OMVYga5L.CIWA@g8B6..PM@-K.;^LK+>J_.f&[I.dMUM:#ZDN;Y0a?cc6
];@0GKZJ:b#WRHE>P=):B<10:3?2R\:fM(U8L1:8C7G=TKTY#^E8g+Xbdbe70IEg
;+H_W-7fa+VMVFM6c:8QU8<15?L0E3QF\=G7WU&(D(KXUE]E>VgYXV_/gG5KG.+R
_VFI#82=MU<8b/d@?55G<gbbPKNOVWCBgMc91D)KUd-6;9EG4N:X)bK_R/06#Ig0
e8W41:Z#Jf]<bJ@/(5U+6;0?8:,?ABBbAS&,bCaS9\03EW[1KR.>@+/KL:IEX>HE
/D/A-P0T+ESXYW6=D-Ve(MT=.(&ZG(LR]]5N;acGS\;f/:&^AV;gFC=7=[B_YL#Y
:3gFU(@MKf0\E2&F6g6eP]S6ARBVQXHKAFR)8?K68ED4<23R]6]OJLV+K<J>;?6C
#PFJ8<V_+.6BO7RcAXKd.6KKCF46N3VTfCB@46ZSZ=^(_;Y==[/Pa70eV72]e><X
aPBN.K^fTUJM#&&IfI-+9UFO;T6aB)HYW,N5_7T#GX=>_U_/5C\?ALSX:A<&GU<g
A;B>FX#@K9WV/NXeHN[dEe.4>2<VX_eAe-ER,/(U1G-c2L6^Z9>DF8Zd4fa<,_=S
.#.U./Y4.U>/EHB,CM3\]X_77F3_2#.@QQ+ASQQD[]U+?Y@##K)2O>2Xf]S)P2\:
K^@T/eMffC99=B-=<BaN)C(5+ad7P<BHDcfX@I#@ba9]<XU/DC#DPe5A:F=WX@WL
CPDS^A5HdAF<AbJe0=Yd8dA-ID]3e)RE^J\:9aT33_SCUHUFSaC3@RY[-6bTGW(Y
De_c)W9.dbf+>CF@IMB9OJ5>KZCH;Mfa)KP/>7JUR4+(Y2INR[bG+N8fI-1[a51F
#=(<M<0+V.XLdYVW^?<?W(9.:;Z);_Cb;R3RH\PP0Q\UYb1P3d[S6C.5S[HI,1eW
SXKZ^I>=;fX2c(L-d3M\6^S4+6:4NfbS\PX-4ba.CS-C26J:GTT6cE]^3[?g#[NX
0&^;W]X>S\;PLP&?MRU<DX^ZT#c,]6:H+U<N\:fOE.TfJ(GB0TR,H2;GWBX.62M>
@A>V8b]ee(R8X4e((+&2HF\N6g_>^+N\f,;E1\J&W1d[^K>fSHKf4FFE9Va;b,>>
&.:EKgDZ75MY5H1A;#==f&?=4ZB>Y10WRD[DL]8]Y>/;H@_b<cLG1TD^+gDde4_C
,8SJH3g7T;BKTYLR7gV0#WI;PZGF.22Z4-b_?Y41ZZI+U/R.NX&(ZA/d@_8;B]+A
>.=4CHVG9,VX/0L<HJ1F/(=_;(9YJ;RIL0F?BRJJ@:I57=W[WX,.:RY&M>7Q<\aA
3cbTIV^9dEAVQFI3:&F0eYg>@^Tg\]c9fc,P^b)(gM/I>L(-eV<[X1F,HSUgNE(T
&E<D8]4eLFI,TY1Pb+f8:J=87GE56Ke(^KQ8BD1S8@_6LC.SUZe]YTBaC7O-Z7S1
PHGB[2Qb8DU)#?We<M)a2/Zb?AIW))8D36+C-]H-RD?0^\^MgdIS,,,+ZaA,52_7
D4C_\6C)N:LDNLT:72BO_Z3aH1L@cV<W_88aA=>L]&#N3V?;:-FfUK_aPcN2G2P1
)X)EeWX(RAg)^<)[7,cgAD?>\B_Z1:TM)Jf[E]M&g_05G[O[)/Q:^7ZND?&<F:d?
6d#XUe7cYV@^=T(>.QdM-].9gDDMRXF&A\FB7cWPN-BfQJ7KI:Bf5TG:DZeJY;W8
<UVJXD]?79<Va:dXQ1#\X&RNUU,BVP?B0WO.4.PL;cN>KW>c#NeT]Bd4CGNc(F^-
S6U&9G>,[8MCT+:&RZdO<P0>^b[&:Sf12?O4WO-4=X\=,HRb^?MgY]J@^];:L6c&
Mb99cN0W_L7e_)G2Y]dfe;;]AcdEPC@H(2a-UA]D5d62EWaT2U(/8=,MB#\1X.<J
4=CEA6)C([Z/&=N08e8\B/L]VZY11N+P8b:\Ja?W)Sc?+g_F6[?X1&5^J^;Dge2c
a(;-)Q]MAN9N92NI#NEFbDV\P0UP5M2@S:/)NB=6c6#f9BW)D&W8<-e\&AY,H7V-
GbTZ91b#3LU0&N-9_Q./DYR9gY<@IE_#-SZA__YWXJada9Lb=5=ZK7PQ\<2g[CZT
75MPf9;6EYd5ZA4D:SZ94X0LWbG2ZV?D.8>G+LB;;eOKK\cBGSb3U]AfSMK_3EH_
Y4ddgCO5SbH);H&EERRa]@:6^-S];8B9IR]-5B=+gf5:faVPP2YO=SR^\MaL-g4H
O#)S:a4bD&bY?P&e:9cRE9BGRCbQX1.7ED5]SOc]g-0O;SNZ1e5L>)BdVNF.[M&[
NE\JL[8#8^8MI=Z8g4Y26fFA7S\H\\Y^aa:Vg.fcDg+_0bKER6:b:TEdNM(HXgY^
7E&OI;PQSd9(R8T[TCM87WGbG@H\(8ES7BNRX):G>E2aODg6d2Z)ZJdAB4Rb)UV-
)F,gMRb1(8C;2[;(eF8QG4V?(c:C^:dK#T7,PA#GYBU_edT+56RKZ5eS0.GI6;V+
\OY/:R,@\]_YdV<:GLR)bE;K3-0)Y#1TBT/Z3+9BV[a4_GXdU4WL0e\J#&4<)N0.
<f]P^/KD&\6ge2P(1fG^Z,EOX+?GO#T,XEb=7He<4#4U3#F.@7)K;Y)g4c;0VcGF
8-8KMf^67/XSb0L>[bYgQ,&;?2GUBde.+)+.?:IBN4ZQ?GZaWeE&NZO<&L)3]>,<
_3IOF+2ScZe8=S4/g,8-(AHIN-3B4)dO3\9K8Z_/J=9M-=d#b9E;I[C4P=;WK[eB
Ba0WGB[^1N2O@R=N6:-BR_B\Q0K:CWD_<XM/:Jaa8d3X/fIL&TcN68Y>TS:eA-ZJ
USGe0H4E@(GV?LB-L-+127gH75Fa04^B[Ecf=@P]W(KNBI)73ILAPWbL6=W2g4@@
?2cOMWL.8gX0;b^)3;J6]=F^&>6AK#CCP6-MF8I>?13DU<P<Z>#,dafNDI&g51V]
:I)HIDF#7Aa3.cL-7:a8K;D2@OA,]7CF\1B[0._A[>_/FL,+g;5D<7[1J#EIG,?9
2A@5Y\Z<Q^7I;Q([UH#98#J8:5FGSG(W[@R#+4P/TXH@b10a]A+Y9W,2+KdMF::K
=[96\#NbJ8X/7<g<WZMB)cL3#QU^5BK6?9Q1-G>,D]Bf>HcM>Z#J@0<DK0)#<Y_D
EV;2f5eOaF/PVVJI@W-CN3d12PV?:F.(e?\_GFg<?)bWST<5)B>>^RD1b[c_+-Ye
&8/7Y#+#T:)&9U.FVBY]5@^[##,4+G8U0/2P9J,K[1CaU)EcJUTYbfQQ\FD+I:8B
K<9IHc5bOQ2>(47NXNZc^5-7T>dVHK,#IH)\R5-[;8@)WR.KdS.T82)N(+0PNM<+
2<J?>cY_I?5d:,O]<FHSKW_]gU)(gK(<5G<(3X0D(gR)/5gZg3@f7A94[CJP_2]g
\1FFJ_)#5HdE_OFCJ?==:Qg^[&4EQbV_@FM(SPRDgFbZ94eI8]R.OB&AaRR89^>S
(e+MLKU&S,T--#P0.PN_\<)(M&8AD@8\-D4)d:;^4:@T)F5cP&]VYS@O/WZ_fS#N
6X[@=/c6Y/fI_QU,>^NGFFW9&&BECLS))[[2G,G-OgFW2[4B853T4Z+LV,P?I&B3
8b?UZ8^gXLA?JEf6LK6ZR7\:AI-Z]W:Y9c-^KZHVWNC:PN_d5>a66g>]G-\[e>.8
5E+aZ\TIT:(D#K\/D&K^Y7D-@a;?.11,780/;+0..9HZ=QJ0Z/#]FF&\K[@>d=M1
GA7)(<H27YMIS?a-&>FM9cdBdIWWg_^[eK1Y0AEI<.ffWOC;&c4KZE]1?YD4XF9>
>_U=dK,)/TCU0[NNFg09G_e\e5cQ)Dc-&KgVWcXN\36.OI6SWI9Z[N2W\V8O-cKT
a3>=@9f)IHNAUFc<7]b92P(5A9VL[G:X>eGV);I=]R:/+)UXIOA21OD2;8[_3e2S
7aA61\Z]1)Nc[1OSZ2\Z@eFA>cdN_W0YJf(&f=W9W-(L,-]c+P]NIf&N]6UH@US1
2BL@Oe5/QH9<L>Jd]>e6.R#]C_>;OgR#IDW?dQ#+/S]IU#T4,.QKN,.V@,)d3#/:
LgY@?C12\D2AFOA>cP3@6-HGbYQ:,O121-7&P&>Y/5N_bf?JXK(XZg:CbgQc=+?5
B<E45T0PW4dMg2<2(9.27F-c7>ALWc]c6^?9Lf_2cNNA\CaF&T8HUHaG^VJ;/,/Y
2b#/91[VCY43gH6UX#cWffc,OgcO0/6[f@:3>\_6S6>X@\^g=EOK2-P.dgCH8D7(
9b<ZDQSM>;277aBJQ>fP?LY?_YT>L)N<[cP>[bW9>OK@WM7LW._]6-G2N<FeQ>2K
C.ZJW\a]8VHPXMge9=F=O30gT2H<(e?f=5;P\?HNW[?-Pd.K#f-4\ag9+#P;e/4<
Cg@#N?Z@IcB:P5)d6_BV2g@7&IKYdbM6g+&R@CY\C@[+:LE9V(/gIPI5Z]=B>(Y=
g1TV7LH9>\GV:AIB8Yc\Y=NDB?RTaUW_(PQKdV=a3[V6?2:\bE(19Tc@Fe#F7]:Y
AL(Z:W#Ud651:#[e(aK3R(SDeaS#/O@6__)O>Y8-AQVe-:&DGXJ+:O2<VFg//B&8
@(N4WAT,,VWFQ3f93.3W38Sf,+e9-aOdC;F70J=DT,HCgaD0F&dFJ[0O@5N5#WPU
G4QW#TKMNE?WfD.OF6QH1C3_9db<&Y>;?HT:d3/FD.6;FLV90XWCI1/P+7IX(d#7
N0/N+(QENSYQTWDDcZVD8_G\?cLE>f/8(T6OXFeK./#N:<P5JaVFa@F&;68H/EL)
fa=#_ZHbNGD8RQE/gb58aO1>R73C<1eNR)5g/X<Q1JW;TE5(:Ng)/IXQaK]=SFO4
C-a;0O45,g1[K:71WBC=KOYAG0L(\)#QK)=R-W+/C19.OUf+a1LVN1^X6/P4]Oe=
M12b3U\,KUD^3KbLE#LX(E:ZTF8FV>Z/bKJ+cFe62/&6SU5U?1gf4RZ8K)_M.88Y
BM=W_dX_TM]fB]g.O]-2<:0&Y2_7I#7P:^4eaA,UeF8;)IAX;HG0#<&JV=Yg^0X,
GR-/Jb+H&7<?LZd#[KL@eY2R?6QY8O:LD/1H_\>L8c=>QG915@?fDa\4Ta[Z;F03
1\H?8YE0HZUfL[#6@G<cDTP;1K)8fL=Pf?@<R6/_Q@bI.@:7#<faZM_B9_<[;M#I
Be39f3_G4M/6(Y2<&\8>_RNGc5H\2g1:]D)#ZCSPAMd7WII+T#9EHO)W[:RMB1RU
7)FB#FW\(cJ(O:UHGD)V4J:R=Z,G&=,/_TEeJU=9Pc;O+N?Fdb#FD.>d=d6b,-:(
WLT0O\1Ze48S0J.<<_S8)P^EBDY[5<#/-EOX3<9Q=d#UFP/YZS@2M58_5U?5RAMT
<cAO#I)^W>^(@2e6([dTOY5YS^fd?WdR8IeZP;WC7Uc:5e7(fM_RLf7Y+II>#4/2
]X:PV(=_)DT]70227/.Y8:C]2;/MZTO-M?O83NW:D\ddNgdS__,62Y=X.RBbK?0V
b-GQU:NPM2W3/71]>BM@/K0UZA;=1O+[MMQX?_5Q?<^]F6g8Mc_gQ\SBa:<N=?fC
Nf2GGN7O&P]8MAE.PAYHL1LAJbHa#0X8\.aTc)SK#N-3R1US7_d9Y#Vf:]QL.>::
.X/Gg4Q.a4_AT\,7YXYD\X,PIJUZ\+BgEB)@C.4@07GK+fb]/R6VP\SCV&\gKJW?
e2I&G8Oc8+LL\2^7U;]N5AGFUE8X+#60RE3T[#UgIAPW3LJ.LR@U(9C?&S/AN736
/-F[Xe[G,KF]+\F7cSc]8VW)-=1VB//VZV,0WFLNRD4CK6>/+KJMHa4fRUd90U4b
XbH\Q(_(UOM=c+2,W:F]eCV?C.\;fL>g77JU9CZ;g])\7eTbE0);XPaFXQ]Z[XKg
NAENH/A)PM>R<1Z5X0\M._0^3KDK.PV;75.6(?]#[)])?C4<XcTbIX&3Xd_XAQ9Y
8[0X(=6cfNX=<e:W+Q7\N05SeUA.HS:SfP+9ab.406U[OHOd20K-1b^e0^Md+=0,
W)0b1)32Y\)cE_K]K6=3->;;.Z?,^_[D@fF9_d_1E.UT,3.P>;g2a.2HSH[>[2CZ
I0Sc,Fb2UG=\LD2SeCeE1e2PJaSX90F1X7S/7<,RK?Mg_W8\-&,W#6+YL,IKT.C0
X3RI7_T28b5Q[.)fe-LD9J/8VE6X5J5CD<BPa[9Ya5;0cSg:D<^W=P0H1<DH;HC:
DOC6JJT&&F5&BQa4T.5[fPgK-(,A+JK_4<Z#=J@HHJe_+O&BIOTE;[5O\H#de,&b
^8B_#\1aS)<7Q23:>^:1A:83d<]EfZNDB,ZJLg_SKM:V193bABBSB^[SVb0?ZK0N
_,?8AD:++O3?KX6g8P/H@?-Q,AS;SZ;bW.?^DR-OdUV:LIEI[R6PaQ3]^2(&\A^-
I^MUS4TbZZE6Y0S\<=P_M<ece&dEaRJJ89dc[B\QU:WIS2a>Z&X:aLR+6#2X;JQ1
<V+TagC&TGB&_cgd:?,7?5A2Gc-JM7;Hd9]2?#UD]<TE4U-cgDW4E&5(a9WIfS\U
dd5W=C08N)DC7[6+];UMdb3^\#Q@2@RCZ<LIfe:E.0.S/Ef(O?]KC:FMSF3:J3??
,TKbX:)G_&[)STIH^=L.6.a&PZ&_IQHQD0NC(/cH,0RbPE.8NTII?b)\]YXTf2:F
J.(B=\TgJJKR5ZcfT:f?O)=C3eBKT_f,.8;627\c)Y,IPJGZ@-<gYc[?)8/c@JXg
CbgBP\>BX7MHPR?/-+7VO_-2WNXNQbZfF2V_5GL[Q:Mcf.aWXNAP&R4JM6/0J0.6
CN?Kd#[dN7&f1):@QRB.e_C]\HEE9+3E)NBY<79BL(P-M9ETbW&Zc?0B_=/8&OT[
O]+V;#Ge]HZ37EMY[\(G7V#-]eP3)4N7c-b+1bSHZ,3QD<f69ffX_@aEgb#<L:Z/
T1/QN=#GP7NNFIfd37W]O0TVF1P6;[)L&=P,eG;aB?:C#)+SA0_Q.6782?9HKA5b
YOF;&I<c<]E4<(bbY-V7[,LB),4&FAE)e>M[g/,;?ZO,EJU5.I3OF9cV?/L+)?0P
I>9T8PSBb\-?YG(J]DFWL+0<bTPA4K=bAMG5JYP<77^W6^-5./YDZB<9T8,>F0H^
X<31&E<-^)L[JLKL_065D9/7L6<I0+E<Eb[N7Dg55)WdZ60G[eGWO(Za8G^0XOcV
86(7MJWeLA^]2g6_UED.f38EX]d]4B35T=1aOLg1a&:WY0WP;&ELOU53Na&fB\d3
?PI^^,W[PWOE+2<:N2VH0FAO&Z(=/:bR7e76T63]ec4S)(N63:]U2ASH=RbO>M-1
7)dA+T;.gF62dg#S@Gc5?AA.\e5Y<YH,G]Gg=V4VF=4(<H>agdMDK8M0^..;N8W5
VbZ:]C/De9:,d]DYP]AgAJO&5<<d,[T-N?8LY86+e[_YX]XZ35VP;-^R]Md5V.\1
@>T))@0JGQCH6.Z]DOH,R\H6FW5IWUE-OP-;\H7GME)TCF@/(2W_]>VK4-R-de^=
&c&CO1_,):GPDNKK/WGeO<E4DOB=a,MTZ#:MY2DTWE]4)T6-Z?,Z.(e](1<dIFeD
N^>WNf]Y89F(NXX<9Va\^ScXFJda<-W_.)77EcWT@X?9.2A1bDO1V14N/XP/=\Nb
/<Wb;eL^IFMU7;c8.KM532/(:G2eB/#FZ_cF.?/#b]eA=UF95H)585HMY_3,,CeY
C+#MZPY:+E^R6O+Qc=5V6FSB6WYF-E74_Ed,eA89gW]9d[d]9N99^S6IL^G[UO9)
U@>8-9#Pe/Vd21GURQ:CJ+3_81):H+GXIS6:S^#E</T\MbL41PVRHg=54CN;3?>B
KYNER?D?#_=LX-.\);0Y6YQG(1/MeQ1TZF)]ZN44CI[FI],7G@cLU7).,gPUP5QL
F<BbE+05YCR.7?&58dYaQ/cT<V+J?-^?+A3A>F[IfAP2fe22-SSXJ=8BV2@9[QZf
R[H?;SfFHZ1(>1(0[I\FQX490K>7Y4SaWg;1?Yf=NF\SI.VdCgEVZ871Le;#2<@4
LJC&-^G)S7eQdW3GDJ-La&\Z)5&/G&e#<0f6bbM:D6(a=?E=Q>F8A=@EP32B1AL/
7f&TMZZ-Q)()YV75V)]8A(@939gI&6^T5CfLbe+J&e09^E0b^=X)a8f&cMR1>B7[
+#2.D]?V(;/W?ET\Q;Y))KXM.M2=MW.[7H09BA^QFE^Nf?H2ed^+DS9f6;YTM#5^
YL8g&F:+K7,@8AJW>MAdN4GKZbff<1,+(ACAFBJHYBV?Dd?5cf)-W[/geaM)7Qb-
GT._&@>9KOHJYeK(C3KIO/;Q\^HeeF_G?5+Ic8Q)f?M=/_=/?&4<&6]3UN+#0gc?
5I\UY,>6\##M]YRg:TPF,X)6<0IE\UdcZQ9?Qc=PWJS>S\2ff:R08YHKVSOaUPfP
#_A\<Be_P2LB@U0Hg33;PFR&(-)J;]S>9cIQ9T3:MUGd3SO>cQ;LK0aLIJ(L)a,]
Z^.>S#McL9.H3]07Gc=)6:GO2QIG<7DOKdgIOTa-eFE0AeLcS5HJ9K/2@^D]UQ(J
DM^(RAM3CBBEM9caZ&IW)b/\QA7#4:8ZB1)2gN3BYSE^g_YYR0]U+0\6+2UXQ6IR
INL7c6gL1CMTa0/fY;4U4&2M-/\deHY^G5,YV4\#g7SBK[.VSFbM.R?DC;B>bDE@
LS-?SQA,N6<gTKLA@SH3LZd/fEB]fT(8&8FA1=D^VATIAL3Y^5)<a7#(JK]NK.L^
1X=WHL.C8:BfX#dgBNFA7FJcUGGZ(L\Ug+67;]CE?U1STBMRONDf/K=TEJ,U:a_#
IP]aI>F+E:>2N(U@e1,ZNPGLJc.G--g-F^>V;U9c8bbOM3V:<RY<gU8fM#N@a::/
8IBSHe#1f?]=5(4_J:/92#&6fgb#9^SQG/E8^X2]CU=BA2@gaXXgRS?Pe@?=cO9[
bLJQcQe6+@LWFZAKEcN,#2Z]/8:9F)d7-??SI(\g6c\3bXWEO2O<IG-Z<WOJC6Nb
)-NUfb2cMK)__LP5;^3G^2LU-:_d\-_N,ARdVgB#P?cKV-Q1F\Z(Kb?E\5OU&6JV
OL.4@MFSEMV3&X=-X);OYDX:#=TG2Kc27[OUd_272>\\\:3.gJNL?_41Vc-0gNN+
_3UCUCRDL<S?R;Mb/bR._5^Ef6EN5)C0?Y9JML^S]AQ:B+1gJYS4,(I\G&,;O_BA
9].)Yf1;gXb4P&1_23@Xf@9AI2CbW\_,[&9Ufcg5@Ng=)GD60EYDTWS]40B&[g,=
?X<2L6&CfH_a.P=b2@B.;J^OdCL_D>@PJ-@)KDfAQG>-FKDcY6=g(aI=;WZ1_d/D
Jc&MM#^/5&8657QcG30G\V0EN9JKJTV=:R2+>GNO?EZAY?UXCgSJbFJ[Y+&3-PP7
5c)dUM[G48]V93VK\T4FP+.He)3P#f]C#]9@d)>VG/]]RUd[dV<=\d5V7A,Red;]
\aeLeDX)P#5UC72D(g&9)J\,#T=b73U&c,-TMW,Y\;H(:T/YIF-166eQ(Ie2bUCg
1#)C0D(<Q]+L:#0PQ:BKNc2-R[X,6bBK/fUA.3Z=EKB/8=7\#f_--166WY2TWC57
KX3TE2__)VG/WGA&5),#Y0=,,0RMQ-J?e0@5Q;:F24#G0cZV(?d/gN3d+Y2W(EJB
80^AYbFLR/4FH598B;/]d<R2_eC)b3[GLGfTS;YARgG[T4X/VTgIWc3#9,C-WMV&
g(O..XP6\J>ZH]L3@DfX8436@a(VQgeT_[F:8__&(XJ_H59F&aC#+9?FLW7:M0A3
I-4FO;g&3GM;+a4N]I(Z4W(gdQ8JfGXC:.P&0ITUKgO55d^EJS5P1\0&IT8P5^dG
LBQC.SXM0Z9S1>]AMg6EfR>FG=+.88=d(dKRAXDCXa7aE?.H4<T77Ve&eEbOQBJN
Y78BA>WaVX2DTc2464aCeIC:F[D]K:=E7B#4>Z]CREDNcE\L.@K;@GG2UKYL=e5=
NCUDa]&(fDW51Y13ML2O9K9d5Y)RHFX)?15N&/N[0A3=>.D[94]I,EG(ET-a?FZ:
A0PYD4g7D[)Pb?BRg\H,bXS9f@;V:/@6fNW129_C_?TUId9.-8;HUf)ZPWe,XK+f
B2e6JSeI@[NT[aJ9A+]\9)\5LdJg/RIK<MV].L7-GTaBO[&.Y-H_Z&]Z9+XO6G@+
)BKaBV9=c((V8^/_>>>7E:>D^[\/I66PCfR=6>bA,8H[6]WD4MTDgJ;-#Z.R,c@L
Y(HFF(KF2d3F9bWQ:.8Y3F_A^7CTdePWD0Lf/#>ecW-;a[<=Z0:EEIeeUbV(I2\S
TY;d=X-0+B@FO)(O_=\:N&729LT#=)7P)])102-eO];eI@ULb0H3<ZC<[R4bf_1S
:5#dc3<K-^;2+3[O8QKTb-LR<OM(=IJ.gQG1V)eeS^B5C/)_3,+TZb^dQ-12?X3O
)Dba1G&b3(2YDOEe/HfJGQUMf7;]<b(;4M/>-A&M;W;^96G^N#:-?Q7Q:)MDHcg,
8[^d:K^TUd7&Tg(?dGS6^]O/Bf:8V[Y/^ZHQ6U).JBbEdC2#/]VIH^2S--(Va+;<
Eb^I(YHPSffL85GR#MF,cPOSKT[OHNB)g#0;F03.B4dHd:R^4[dX4I;1cW0A9\ZQ
=7e;gGT9ZZ,L#d4:c.g))>:S_E^GK:MfN0?-KG<T.=/-A/4<)KWBDFWPb_@\B5WB
8Q<=2-PST;2>1ZdFDf>@F<7g_UL@>^.g5NQe0c(1#AaaM>MJE1QM(XSF^HC(PY2X
Zf]KR8N?/5QN[^A\STI<)DHg]5R7(RA,RXI4L@&^<;@e2#DS2I[7QP2?=L@Z]a#f
L?>gL)FTdgE3;HEKO>WbJ_eBPc,\e#93]44-d;<Q35=59F:b1=a.gX)W:5QEdOeW
R7E[F2Z7g?WIg<cM01XV]L&R7T]:&AbCf]d+TCEHU\1b\+6&Q)(e;[6bRKI-BIW7
J/Q>?.22GX-T3_OGO4G34aU4>KU=X,QW5c,K).Y-PPXb#cX9H8(PKWTQ?Y>^]^gc
#,\3,,R0+7L(R2F(_95UCb=3?W+^_VIKJZeAG8MGY-e;NWJ\1UC-^,D?P,L9Q89C
-,XO&^XC)<03ZHX[>_TL5G]QRWI\(g4/KTDf?;?Pf:U.9dD@R,=6-60W=OJ\\FG7
1=:d+5PJ_7S;cZ3(9+XUZ0@DJ_A7#>S1S9)e8PWE/cHQKK6_L(/0g[0_>,7QBA9>
2HB605#>eN-)GF+0e,5-RHf1KUC[(\>?P):KVE3_^._^Pb(:6E_SRJGPOYQ5B03g
I>Q9R&@Q><bcD#BF:IcLX@-Y0B?.bDd9UDf./Gg?5IJ@QJHg#WSMVRP^.d]a5VeU
/\1\WaB5MP/eS3[B[2gNS81d;M;e9W]EF=fO,f@M7G>9V^,3]^-gaP0.S&EH_X9#
2ff.TD)[+8UA#I,W5\[?VWbeT3679=\&T+W6<1(^FF,K69Qe9_0WV0+<U5+Oa7PH
SPT4Q7AbV2(3GN1_46(,/WFP7K_d)+<KQg8c6->OQgJG,1&,V8Q4]^IK#IG)RcOd
\DH69UZ\J(,Y<VH1Y]gG2,MU#6O#+A9L6)YOb;K_Jf^BaTI(235K2G.YO^1c#3?G
G#ZcI-KRM4LP/Pa-HC7I#X&QBaEb3@_L+++e]G-2L\G([RC>Y=@+36H233O(5/2W
DJ.D>3791Cbd+>0DRWb]VI(eL+Q+Z0SMa(?NLQ9XIEDB^V/[P#0I\^#-cOb;#\5d
([2g^C5[Se^F@QQ)YB?b\(CDWTCN2S7&&Q8@PBESSB4/7,K0fNe-,/99GZL+W<&6
a=4]K\gC4)&ZaI#R^Vb245);-dPJ3MP?+R0TI)-Oe.fNb&SD3T)U(P.B_F>_(\@&
]F/OSN8(&UZDOWe7+4#VM/CI\0dgME9Of5ARc\<Tf2gL+?/3;1+V?(IS+0N]99^(
g?4Z@[\<;]Qdd4/UEM4@M\1)^?@<&<(&>9]REGE&#@EccCX=9-ZE2]X4P;NYPT@5
^TS?6gd1U\]=)H_dAXPLBM7X)CJGB2A.5@YF-7cP^ZF<(CPTeL:AX8;C[?TPJ:)(
2&T5eQb1YQUUP^4+AR#a8)HN0UVNG8ac,=[GU=aB(DP9V+ca;PPR4,-&WaJXDBCY
;FgN&KC4Ze^9L,_dea9Qbg@)Z0XHOd#_]@)?7OO1?SV#PG>8B?c,MaL:JGfSQ3-;
J7E<[((G8_89O.=2B0aXJJ8BHC\3_CT]QJF)E[/C_O=A(CT8CBXZ&M&fY33>^aXK
@X3+FVNG1_J8MP_:Q[?)DC/SYH9#]SRGW]5e-I>>e-\19M[TP9/@\GDbb^V]8Y?#
Nf_LdXeOSRfK,[X5[0DV1+_=c3U]Z^D)599XAHC?V]Ea:;\H^<2C:2gJ#-R]b=DO
5EPYKYO<L.9;.5[MB29aZS>7a<.ZcW\[=^UQc5b]Lc_dMP192DH8cd4O:/(QO6&9
dLK#>,]T]acJ/(YZ;F;,BI;#FIAAK1&6[ZJEfZB3TZQC:KX?EZQS+a<79S,6+&EW
72IDLE4@e@Df:T+2I.d-/SYG:^536UBB@G6B6+CBHW4K[#Q,Q[<^2__I(<DE]IH(
fJCJ.3HcXf:X/?/KGGc9F5FALJ[@,?VI7+<P&YEFLU,.Mc5CPZVRacHJc.T1_B(1
<>2]I#Na9X4ROcYT]:8]1MfeU^#RTA[HNDVLQT+,?D;ZT@L]c,2e/CDLe(N41=cK
cVb,BJVQ>[R8SOC)g1GBaaY<_Y3\,@.9fBYH6^4EJEH/EX;^6,5J3RJ&gCA-V7L5
7&RV5Y>gX85R>\)S>S&9.G</#Od[[@?C6cJQ][E2N,MOgd7PJLS\[=G4BBQGX\L5
X(:1BGBR;AHaT(Y6V([R-9V:PB)5Y&@-cSNCCWY=cWM343b^[gQ]V[b.I&1UK.Tg
4NM>(L^D=&dH@-_aT,^cG@CJM]5M]A^4U?P:[CB^6@F_QaSIVdQXZfIG=;=\X@dD
1T_dBI-678U6Z/1PV.DBJb\aN@6>J@L1HU[6-)MPR,3IW_ZM1;?bZY)./a&5(:UZ
<C6E\_:2BMPDV//GCMeE,,T:[]#/C?Rf<<3]eT01BE<f-/e8IRZY>SP,a#=(ZQAJ
:(X&;TG1(_bUXL+))d=VJZA7;dX)/ML^8U)<NM81JNI)a_OO(?(fNV&U+P35D4))
(LPS]R6AMd]eXd\a@AB&=(@Fb<WHVAEf,9)#\(Yg8FF/^aM4B54;#2PKG,?eG_6O
Yb.0N:QTOYT4e\#T/6382b+HB[PXL4/NW@H@;J-DdBX0JVeNeSdHHVOMF=N<LD3I
d.B1+_10d?H.TCR.WB-Pg53\Kb7QP4)7R@M._DAJ=Z0gO7R[^3:e3fAN3@;eA-E?
J)>HKC1GgBU=SXH1a<^gXLab@@2HcXMV:M=@T1dT>g,)?BW?8:.9Rc7-G@:1+J6(
+7d-W&-K])-dGHVY0DM&Ob+NGcV=CY4F4.<JN<-db->^M/.E(9DBW8=P5gSIUSRR
UJ9XO\(\FgVVP#]V@Ug\G;<@FbH&bS/cUO4[-2G(6(A/0S]S<TH]1QTdaR<U1DVG
;2@:D#bcT<97e83].YQDb[RRYKBX,XRDGGYQ4&MC(b,S3QT+d_ea@@(Y=0HaPW5F
7G3=>>M:&]05WSRG+D3YZ4DYG+Ke)bDQ>F5,/O5-/K+5>Y([GH7)MG69e0Qb]5NW
[LR/Ng9;HA7=7<_I<.Wg]<PQfZK#Xc+&7R=7M2\baC54,5eRREWg/TPFe:P.8N/]
ST_CF2K;fDQ#Q#FLJ>5^<9G8B6>:[[W0X8=]S7cCIfdd]T-P9R&(X7BU1SPT=94-
Ba3V/KSc6KE/+\>]9^?UG4(UEPOeM=[b1bSUQW3,@afJLIR-g:&1#=P7f3;Q7Hg9
;6DXfXAKT9gfLKHTga._bERR.<#@G5:@[U<gER8-D(L<b;ca\ZO\UYeU-</ZeS6#
WaGbd:82(+VZ/ZI7VB=]NVAQ;-Vf.19O;Ic6K^7EBY,U74+38-.g<#37RV5.IF2_
3&#2-S)4HE9M<>]QYB-WH_[.+<T3=#EEaMTY9/;?HD)PKWGN>VM_aRFJVc;&-=OM
UUcTfUSXTC+S/PcaXE6fFNeO+g?(3Q:&,V+V5_F[/SBUYTY8&.RXY-X:DI:B7gWa
MMb,N;/AgdN;Nb[@TUOBf[4d@I:09HX8==<M)R;5WD<IM\P&EFe57#[?K@Ie_TE(
VX\e?FLS,TB;L<J230B7=.J7R9Ob2Y.50^#GF@M.e6A,3O;G)=1+@UR=4NT,:@^F
YaQ;]_#T3E1K9?I>dZU#?gYX31O\A./>UQ/eY<Cgaba/GO2P](eM-)Y@CT,_:C:f
N31d_-ZD@/1,NNY32FCM.G0]W^,_+6<I7H,HUb\1aY2DE&(A0f+2)6>=7M5OZ2Dg
\&FZ,1d@GXZZV[c;cFeb0WH[MFgX;5Ra(9Ibc7HV_V9GYK6T-]f3[_e6H;<7QA:W
PS:c.)#CP<;A36gJZ.-)Lgg3A48BWJCcRJdH#L\f&2cSc0>f=PIa05R@U,;^McY5
LIW[f@&-.QUTS@A-+EF5>D8DVO\SY3bI+49=\JA-+D#ZT9=1E(NL\[U^^XX15)I7
ee#aWE4J32bFD=ZUf&XS:LOE)]9Kfa;(3a7B[LTE;ESDKGf,FX^65K+PA@cD&GY]
&N7UF-#gW=(B5d3)Jf7/@Wg>S&aQAU>J[gM=H(PB^4TW_b24_4)Y-CBYB>:V#Q6Q
P_KIMR4U?cC&LXH.LK(8\T;Re;,TZE,2UH>2c20&?1J;4:S)0J2+eHC<U7Xe&1AK
P[-Z0eg2&-9O5YK)EBd,.\)+K(R(#aH6V3AKH,L/+/@W-a<?CD_)D#@_JAaX9HX#
b]PX?(O2ecdf6E-7;;g&>CLQYVSK(d9&S3_K]Kfc4E4#?0eX\\>NTSW0e_=^@T&/
QX-)YE&a&1L&1\1caZ@C0O(,HbLf7X_6Y[WL0,Ac>S?]VDQBPP\NODFN)7M@gd-I
NHM/Qb&&0[a1PgF+2+V@X?)f1:?1ZK>#,B:9-178gW6SNH[Q\_622:b8?6D4WAcf
T>CY3DETb>8SN:?[JK4&fdC>:9=Y/c1#d6H?CFC]OLcX3_@6A;HY:6Yg=W>38c66
1Y1,E_P12J\3+L3Q5BJaLe/\Nd8eHT)W\7^.N4/Y@_9G<&&2fbYbgS3bQ]=7)D=+
OFL+K#PeQAdUT@fRB4+gK7B\)Q[,\SOCQ[@\L+.3d/:J93eWXK:4+g4FI^56?M/g
,5U:f?42O,X?EX;KP_,E8/VQTC)\_;R=eZ@-\?A&cbH(NfI4Bg[VZC7H0CSf++O)
)DK72=5LG=#EA/4RfYGVZ&=OHIX13?VNQddAAJBUA1>C?QAQO:69[_eE4D]WMTD6
A,47,07Bb(cD=1-03Ke?,a5f7<b1D;5c6DN];V4.R3SHAUZ^&6O-cXB;<X#()]e+
T^9DL:GgH>^>cZ-Rg59;1:(IX(TDT:21_8)^[^H6<L,d8dVAQ547<\GIBGS(>F5a
7(YRNbKB7[>e-^1OF1bRaJI-ADCBYE3e)g2QRP,\,04#N8_BacPZWT?WZP&fc<a5
KOG9]b]/d<K#\AZ/Gb<Fc-82:C]XaY8K&cJ@NC+[K00>,KK1MNA5/1]c/)e)8=@d
EG2Ye[8aKdB26g\F&(EZ)0O<IT;=f-Hc6N:)8]3QE+ebXCAf152gXDTRPcW2PC+e
-[A7P7ZA-V=G4Y(EQISC_I#0;=WK-#CJ(Q7eI&C4KL)QV^W\KG7?@N87SJK=^5(:
8E\.K#?g#2O5\+P00ZGXHI_g[E<02XL[^A@4-[G11/MFd>6J>G[GOC.4QGUYB7Ra
U38c->W,#?7<.C5G1[I(+FeV_YbdNHa.@;U^]YH8=adOF,+SXBIQIO,>8@&1UVLB
d7ZE(2cA:XCcSgU77<.:V;afJ^Y:Ia=8aUaZM[_Y@:FK4,+<N/:^_:85DVadZTU9
F0(+23fPC<1gI=UPMB6g2S[JcXVV^73R\VA6/D([?SXV]#e,9_<>1V.)PNLD8J5^
29BMV@D?08?ZY4-_b#/fGgHQ5bLVC0#Yg_(C#N<BEI=?(J#eJZbfZV.ZOQZ./FT(
K](K1^@&_X8Z)TMCEG<_CRfeg&_gYgYP0>.);dSd5]H_[DFA^M7AgegSCd:e:d[N
NZBBTaLSMCFU1_&L80b0FdNM_A^CP/1CYW.-]>deO_ecBE#K[O<FVI+/VUG]b&3@
?VO]---<C-LJ?VWdbBKV2O]gBH,N(Gf0,.[#QQg[#8N9W(Gd40dbM?LQ1M4/a@;9
81MIXY+UO&gB(0D^Y,FUJ3AX3?3RAC18?B9e5Deb0/g@_>)P+QR3+(KBEN7Ve#@&
AKK60>\H=M[>U:7._\75ZcE3B(Vfc3N7@BI7=<@<2PI2(P_e9C/AFL4NXa9Z(+1<
56VOS8fZAJCL2A<D.X,VfLOIB1IR&:OQ7V+[AdAKXVT^C#_?fb-E;DaX9#:H?A,V
T90[DVKH:>@CALO5^VR&GXN6UR]\?d13)+(E?dT]PAC;F<Z4c,>47ZM?.C5_=C3F
e98YT^R5D6Jg:f<V58+#)fA]ZMaZA/><>UZbGKUD5Q4M,IgdGXDK[&Q5]J@FV40S
dE:,b,=@e.TJa(6,_Gec>8=#/PZ\\&#3.Yb:+JE;5_Y(23RT+A/MC)(#?)O-ED4L
WCAQN)8A9TaVC-&LH5K3.37S#dV>cFaP1Z65N=994<b-ReHL_/P[?,Ab[D50f9_<
SQI-D+V<a\PFaYJ7?IgGZ@M1WPQO/0(&/W(L<&TJ;+BWR8UBd+-f7J3?:8Nf<3Ad
<S_^[I](Y9A97WY94Yb67bdH3J/147/&Lg<ZZC/B3Z7:@:Sa_1b/17]FS.gZ^?Ra
EW=[abOCEN)P<M3WP_/<c=CW@EXbL7#;ca1=\eaQ\5FALNZa64ET7+&M@K]ZI,f4
(>8_=KdC][W0\=T.@=OeX5e.+(8USSI+1U^3<bKP[XQ)W<5^(HVXf#8H)BU=,T?+
cdZ2=cWF9H6b77=L;G7H44Pe;]H7VC)T3)9U>:f+CPVXMXOd=VG8-+cf(AP];7IP
3ZK#>>,O-9J_<N:4R@+W0\P]S:DY)eWRd<7EV4BE?,IZagMUa]a0\6E/H4J(d,VO
Z>fRK6R\H7;D4RNO:Z>QBNV]#WC>J[7H=cWIfSW)J7a,/@fTe6bFYa9\.5AWCP+F
g8#1;<)(39@6]J9V87K0CVQD4VGHeP-Z#b.+)9g]B?[EN#bYXZ[XceQ1gVD9-HaR
?g0=?dUS,1DIXA#)+UI@<LD>Z7c-Y0:W#KL^_+HJgB_4Z.5#[20BX[UM8-/UU7a>
/bD4&T6IN?B</IS3SUb&.->2\H.46><KN=V)AV6>^,<.2Z:\:Y:)(182a,@[M79N
AL]<[[2/I,,]2?..&GE?N-cdW4Ec^?9EKRBJ,O[8Q+FfT@SMI\1eS^A=16aGaIYO
]>ZPD0#5HFX8-&d?62A3Jd7[5N2V:>3I/9BBST.577HE3T4#J&c&Cf,57L]S5+^Z
/G-BM+L(3H-?Te.5]]1Z&dR\SDE)?W3N;.VZf^576S_2M]BFP5->c(FH33=&1S@3
7,0eC5FEL[&CE[EI(C6XIeAeXP]<5a-JCZUCS>3S1]LbJQ=SQ^I(LTSC824Eg)_U
+Y?XHDUGM4E18BdQU_dV^-=T<9bBgRZg_X]2FMc2)Dd85L0[b&UG\CSc>8N2;ET]
g\M0&/#7:CW)WX^.X)-#9-B;ZZ-c;MSTCHb+QeR\_VZ&YPgb[A>6-JKN[7V9X.3[
F@&51#9_OP)Z4)>C2:SdAKQGG\^A+Q0M,:BT_I,M:XbC.Q@WIeO+gZQ+b<g^#EQ:
^GKDI>=Kea;UXPEcT.Te;6d=2E825e;+T,]#fCN?EDX4_Z5+^QML)5Kc#0,P)F,@
@)F9b=gWD60L^004W,GR6e7Aa7(cW.W./YI#NNY[@f).><:De+-?NY?J@@/gXSMB
fP40MIR.4/Q.QZg_:50=E8DDcVB8GTFOa(M+La)MA_c+R2NALII8-5=NWBHJMM[9
.73+eK\?V]eQY@J>M[&Y#M&\U.&Y>Gf7b+8;Ec-5KRg^PP.g73J_].?2Me;CCL,S
VPe,0BM,8(]QDTVG41F>a#9.4)P?g)H&-UXX<fNJD3O.69Pc)[cALY6]J9?>e6[:
,LO8W)Y&8.+.HS1Wd_E_dQ^C[XRW4DP5BMN&2e1<d+>:Bdc@(04C.,bH(g]K63@f
7]VfDcKR\Y^,GOfYGI/Q]1EZ@Lf7SJO,IZ:&6XURFe?-_=W\PXbAJU4[=&dAZD?4
R3A>c>Yf,eR?=V)bbHgCcY&-g688G,>,(-WPb5\+PQ)+LD5LZ.\PdSE_2H.BGCK^
8F\:O[;Te+D#/f:SL9O)e)O9IPHL\.eWY4=?;GJ#?[8[dJ]IZ(S+)VTG4LTNbcF+
L0_dH6#eJ3(Q=:HaMSXK-b=N@X(<Y,9UW>/JRUaF[(;(OAd[Xe,6,XYZ1I,>/(]B
aY2)f9+VWUV?/>BI6>BP:NH]BZ6]I/DV7:KX[7&5FV0;g,4BHOgeWX_eUE5RUc^(
61=U0:;.YK?/DXS(L4Z2H4C02&Z]c3Ze@[;GR2Q\0?Rd==?OZ)XWZGT/4+DH=AE(
&e6;CZV/7C<?QP,gK)g^]ANLQF(2\@V\,6I9g]2&>gY_ZSRa6KD+N]16R1]X3fVA
X1J(M&57gP@1[(9=40XV@CHA]>VU6IW;ObWG=H_Q6&.CYUJ-dONB)IWHFRb.=.a6
[;.5;L4HfY/ObZ=/H?;^@8CRB1E]PF?JH1[=6VZK_YH:?[&VHAWW0:[UeIPba3;Y
cKS\&dTRfAFA@(2.b=4,K=Cb^@(SgFVVMMCQ+YPdQICcg)/>R<R1N&JK9d3c]Z:B
M>7@,QT/KdGK0O&R5Df?B_GFg.AYaVL>+0V.M^bNY\)2Cdc6QTBgF-B_VNQ+d\(&
WGCg/HX9MWA9QDE79a7HWeRG6+GN\b8K3#VN^-C.4&NEf2^+&M30,D)RIg)C_(Jg
_5g43W#FQ\\[5(L0R5QI(83A9KO&2C[e4Ib]g9-KC0fR&G/eS)_aPJ5)K/S<0:#(
/RE;[g?=eA+/Bc,]&F-VXL8[/U-;,S\3aIY\-;6IcI9_c:f5B7>Fe/05121)95EP
.5e:5[SZ\?)CJ,?P4?]+;3&YP;aQ[@AC-3[CF_2YVM,KL=:WI@g33@@gTVEb3+@E
[)eF@#BHGYe7>gP7L;DLgF9aJF0-.9[7;]8b^+[_7I>aTDX)\Y(KUF+77cHY-M\,
a]+;9IEZVO<5#AfSWO\a/ONUXQMd4FYgW/?;/.&RX.-::Z.7_LWaVQ7L@e(^N&6g
=gD6[Kf16d9JCJ)3)g.@IA0,Q[ca]QC6b]\F&C/a5]1;Qf7XB7ZS4&-ERdAYK)RQ
N)3-QO&JZ0#HMWHC2?T<FW)BE;7e8#MIR115>NM+bdec?]cGI/?8a/eB\ZWD<R.b
VH?MP(T&:<Lc@8f3<QO>/:#]?PSY,U1_M<g>Y0-128>:eK-7c=W>>\<e08@CA/MZ
;8)UZ_+U)CJf67W0=)40?T;899,N?UFgd2@,-0DGBA-LN2f)SgAXC(bULL]/:]Z0
0/Og&-dZdU6X3Y76L\@Wf,9FX3SCWSY=M^XE2+4FT8S&;7@\EJ3QRRV];Ug);)Bf
3/:Q>0R>J4^)#5/0325\ZN:FZ3&7b++P81J8RcC:1.4@03][Cd<II&S6006)b\&b
?O<9(CU8F[FKaQ,07cgf0_=TH9IBOC?7H,&TYO77N.8D@BHF_Za-/GcJE9FKV6Zc
(gcW42SZU=KP560P6DT-VJeV/CX>#>^TGD+>aLP.Z;g+]<A4LeNg)9G7B>Z:;VQJ
9cPE(8KR8eU#/HgHN](YI/XV<W[XQYA@+:+:(CeJJL1/X\TOUIFLN<N)[.Jd9V1.
e??-)e-N)NM7E)-4SC\XD@b4<1B]S01A?^ESba0EHc=([MSBb;OAe@##4^;#)ZS0
TaW&5QGMe1?;JI99cIBDVA-OC.,3g)^:?)#2LP0(.gcN(+gV?L()[G2W@.S&/1b=
21X2CNFG&;ggEd3X0I(O6VNOC-AbZ;ZLZYS.PA],R./^=KMG&#0W0J-E7\R5>NQb
X9.]5eZc-6F([^+_&=L(L,&bJ><&IJ2N1EO&<K0/YLRL/)D^TE+b^P\[Wg:M:cMX
Q)QQ@GF48B^_^PcXfA4,WNB#<bAS4e:AbYBe5eVKMU[F]aW?5><\HE.5W8;W49^N
QE(O\8E0;4/+H@D[bRHR;)>.-YNLSONCZ&LN_SaG;T?)U^/_>=ZM0@M8Ja]DDPW9
JBA>^,370gP&6JMObW?EINZB#Mb.81QYfa5,QD>\fOI8Fd_=ea;a@b3V,5a-LG=F
<[0R3]R1&IN(F69@eR\cK9(SC^6bP+F[2)HD,EQF7#^4\\XR?+5K8H=?Y=T[H>_M
N;ga?8GX0-==?9F@e&H?2HWT.YIB8<Z&a8LZ1_^_UNT>5Y,4:/WE55>HFcV@])MV
.7P88BK4]-#AW\;ag+CK<AV9X#fGBO=O]N(-WJX];>9JN/8V7eS3S8;TR)R=e5A(
>:K<CZc)fcZOf-^NO&g8U:gdb]VdUB(1gR9B;#3.c>GZ0ACfc38RbEK>d#fXC1ge
(,+aCL<M>LD2bUC@77@0CMRUa<.(-=5:MYJ-@)e+8F@P_K[63EY&DFF6/&dcN7Wf
\+f?9K>2MZ[_:UM>c&7KI3bA29geg8J@FGV+?S3gUYT+.bR9+?LGCP.)S,HfJb:&
H-Q4Jg@<]\^\gN37RV8[47GR<-W\A+^PPO,f8W@B<5dN2_e8K#Q2U#b+?g22H5XK
ae(Y,UANe=ea/;bBM1aR7I9Y^H3,.NbYA2^KRdHK4S732/>&S>;FC8)0Z6F_-/S+
19FZ35@aYId15g@;[a+#^ZGBV(OD#TRY<7LSeR)>@<.[+-,PU+ZGM-4^XYOJIK;V
aQ)3P8CNf@T9=]>FHeOD_2c#M[F;2)VPF2e.E]/_[RMDWXI;:+[KFZ7g\8FXf9H.
PS7=cY078]O4&QP&K2T?>]PEKFQE^PI@d5TUZE],1(g98A@0CC\M0LH5=D:Y&VX0
<IW?_K-Ed;XbF;CBP<OGA+T<1MOE(d3_^T?3KLaWa/7]^5a8>dU4Y5Z.LM25B9;+
3cf>/g+I#6QD4c/J4?/K;K]aXKI&O^^</d0V/FQW>J8+-/>EG]F5V3+=^Z.]GHOK
OeD+6J@&1S4Xc,933L=LSLS>W(bR2KPW3_1S#MSP4F\TO7[+\bXST8/,5&bX0BG4
?HeQ\,I7+AJI+Pb[;^\GT.8V5cHY(7,^,b]\K&4DaAK:A>fcJ)CZZf>&B;/DJ7_f
/,NbC@+I+d<a07MSgC^GW^,0@5CZ4W<ITI&O[QFOaAN6aYA+e&UEPN([EZ(/AGg]
>KH;_RP)^24DZY2SaZ,XS9NX8\GYJ&5LKI\@:(RJ-)L8D+S8(I30X?.A?)XX=,SU
&7@4)B#<O39V:=0>RJSUK\G_J/f__KMIQP?5Sf#+<CB5Wg9R)O<E=267RSJRACJg
(e9YQBR)O23&FT#dK7fG]Y8S/XQ@b0e@UU(cSEU/:3VGS;RgG7?f)_bJ?ANRD_MJ
]<W,];XA.=:D,V;3>dc1^SLb5ABW3NVH->XM#45=9-G3,fW48QCaRTIHXMSEQTOC
a7D9@cJ3b<F=PEfdYWb7,B,<5+/F>V2>M[]:RAJ;H)M6G#I9)acbd)USC>DXH<Y+
TN6J625Pce?7>X5@KKR6(SASLZ1dJUSMO;^@C\aA6X/-18HJ@5SW09J0:JHTV#\M
OQ3)IKFf1Z,a,8WN4L\^QG@Z^;C2E.c@UA<[.eGJe0^F9S9TE#BRK(W)-#]g7DK>
g)B^GTDI==_A4U=5#[+4_e=.6>0B0TN(FfVL,BS9:5LbTU?=G2/fB:#&_H5REX[:
-TV?+f5K,gV]4PRa\^e(X5J-QJ;VVXXAGH;GY?2_YU:-/8F6,EC-Y]X<gQ<KW;Ag
.cMBWZ=+IV5.DI/g9T:L^Ha#Tf5<6/G?[P+Z9d7e:RGG0P;1@WcG5&8>3+b[NTX)
./OLcfWX7/GI_&A7\(7X\+U:325W-Y&cBM#Ad/^K463g(a[d-b0V;TJC(Jgc_E4C
D[Y?gYN+c<Y;8M.8O[DcJ(GTOKN5RQF6b1:/O<Xbd\6L4+(<LFN@cB(=1KXB/?[1
@.+@L?NCX8MTd2XD^8=2<+OSIdMe3(#eCE:b(LGBM>[A4_>#+BVgEG-@g.5\<Z-<
d6cBS\W>/eg,8Z)eH;Z2(5B(&UBY#?).XP1@7[TSMaf<PIKcPJ00KQY\gSa+M4dN
U1IO&^A./B0U<1AA,Z>@.0WSfW:4QO(&96c.)&I6#;\K8VKL@-;R@>ZY+03+1BTC
bHR[5@J(fS[:?0W+PR+N(e6(CC[HGSD/#RaQ\#PfaC]+;;MU;P_#ZE4ZWNYZ7>UY
Q45_bcfYQgS&O>HW[Q<P^d[^c<Yc;6,W)dOI17BaDPg-8Z+B-5a_Gd.TS29aG0P2
ecYU2M[YJ&aZP^8cO2OW#0#d_X@>[O/bN[<^UN9G-<5)5c^CC_@Q>8cC+YL>5S>#
>(<^L::04GfCS(K()GfEZ>&R]9T&W@S&6UXe6BF_-6TK&Og<</5TV4QMAWc-6H.H
9VY=51+;N;9&_)b0#a(#d=Ka/;27.8Yf)1[d;.&]:;VPFSN5>=-#ERb7J_.,2?1?
K:aG3R=&MXeZKD>Uf:PgAE;3?_2=GW_gO.+#f<[D,U/B+E94_3@JIZ;<GYdbd)S+
C(Q.Ve?RG,.e^IZ8:13TSZ(d-.dSN::45\\]f#:8?X4AfMH5_?L#/7(>5],5?4]G
Q3fXW8JF\/3Z&L[^7IEaTSK<?)f@;;a/C&Q_BE\P&@,9#:L]G(F;@XQ[^O=57M0b
V1?#7Tg0=H]WN@N903HPa_cTB4P([QKQD]J+Kb)\Xba(>#f>b@Z_Yd9)>FZ3D3J>
5eCgEVJXcf:R#]DP+^WM^Z\+4cS@CEYG]=\CGT2@(Gc,N?]6cWW)2[6CfeC3dQTJ
PFR:gKL8GRQ]3c;)\>_9)^d]bCWZN#UEY,O<O4;_#FB2A[C1NAZB1A&KNVOfD236
cZ@PF#,D(^ag3C8YV7BY3KB\6F=95A4NcW5eQ)T\54M:GJ7g?&fZ>ZV->De:L[2N
R(g,V0T35aR@-WLf9JVR]\5gCg8^-1;:7TJ+_^5a,&Ja.#)\\CCZEa0S2._LS,<.
ffAE,7WGbVb:>f0Z0XEU/f]7bcCI8QFY&B.Y^KB;V?dWFc.b31+EI7[M^;G_Kc0D
<5YPYGM[3-C5<A)G17bgUK0Jf)ZLRST9;S1TaSZfT@)a)1TcF@^_CC[1e6@T7?a1
0IBf(fU/U09UKH,9FNeTdVA7,+HX:4TbAX,9FY.@3)V;J.(,\N9RF-RE(H75<=MO
1GZXf.ZVXXHdR.J&6]K3TF<)6?I7SOB(+A/O2T^fb>-Da,(@IFa5K#6A>:W1S,-(
JWVN6>OPB7UN;-0H/.aRB9_4g5CU?f>#]bHVOHdXXBVY9;0VGS_(P5VV0X5Z11Ye
0-fE]9]a#6a.89(QT8K,FC-[c][4/&9+>EBC]BeSR)-(MSB+7&?A;)M@U7D3OTEX
_<)9MF^aCdb5>cR#IGUCS9Rg80/((:=E3L/U]cKF;M,d2W6Gbd0a=V8ETCRA6LWg
D?bc[C_FT)0[=#<RBe?dQaL<.fA?_BYNc+:aWVU/CM+^Xb3C.-B#OVF-]9GDZPS_
)gBaFVGGMXNAA-Fa\.YGC+7(C7MG5.^cWYLRRNY&27ee5EXW:YEcfZ<+EJSM+W7g
052+,MHX(HDJ^LZe+>_D1b-3A[4#VI^c5@7?@@_AI3IHTd0bH2>.1B&258NLXe,K
OgFeO>8-L_#CI2adDPKaE5BN,:ZG[ScUU\=+e@F6[)LI&SIbUV:f?9\eZDEb3UMU
H/&;aC._1bSWS;3;_[+9H&34(K8]1N]]&GNH6/B:>/WBG[c8>M)a54U;_)/5V:Eb
,KL>4dcG>>8gNXcg?f&DY2HPBE]@C?TUde[6T^A:VD1FR=LgQ5@_da@eHI)1d_SK
D^LR2KgP5YAE=K-NJ,J]2_-#V^5)d+NID=/:aS@@?JNOA[1WdAO=VVc4DSIL[Xgb
bNb;#.0<I7^b<?+FP=RA@7VQaPBR2C#6+#PWK)T2R/]:=L.+1eb#4.A_L+faeHC6
OAIaJHe1gH.1F/=W;f#WU\B?c(9-/JI#5O=Ae@BaNId8/,ZGM4(XdFAc:dPYCOE]
R_-4TcO)8>Wd#VVcTB=D[]@-&6P;+4D#4-C^U5#QQDg]Gd6/L\J))41(M4Z5Yd:U
#9467QcE@O[D;[FI0W34)X]fDT(T:0SUKOOe9:T&+KIb5W+:^^_5QEEg58>_Y.^U
O[cCW(cD7d1K^>51gE(VOcg[)&HcZMJ7>&;XaQbA9S9a/0S]AU/a5K4RLI@D)-EQ
&0QSTULI@CLUK&)[6+GV7dTY2WcB-dIVA_#BVR0[-T/T2a;g0HT\Z27S.,1=014J
6ZGN^#DMN]0DCB;beccNd([P(^^gPGd/N,?5WA0>(H&e[=O_T7N[Y;F\5_8QcDV#
H_ZZ0:bAWY:0OR=0RdRLOSN8@LP[g/P+4NH=+UCKe]-FcQOM/:5f@8TURA;UC6P,
GFCdEb<I>0.8?f&Q@8]<8A45cKMf^ePLX[U_08P]UgEEPOTZO&-[TE&F49d21d13
6M]FJGIaAH:]g>-2P1WfX<]JQ&<N.dQ/YZLT\2F[:\C<,JYR7]X_V=W:b&c1VK0F
F8_47(<JaVKEC(Cb&5525#(68G),E)-EA@U[H5S-A^<S&]Q>d1c3R^D4]@X8VZV2
Mg5#aO5K;U>afV1YX/96M,\)O[S8@S5??6SO\cC[0-fegULCVT;Neg\<+DN,S<gW
S6E<&,Yf2EIL#DFW\JT)-D]21Z\214-\S#ecIE9&CTe,M<D&6#._bN94:c)gg1O]
X)JKZ&3)A/Ba@:?+d2XCe^\O5VVbSFO2^bMVGbAcf&M/?1/8[C\Y3S;?<^V<(U3,
<_DTB._G8];\_]YTG(W)gASN4Sd3eJV+R4.;)R[\U;)5I5IfQ&=(=UNM9Rc^=;#;
._Q<Z<(aU5N,NO59S+AJ^6J_<8bX<J;^cJQOQ)@>=K,-cS?W+O4SICEU@DZ[0<bg
U3U=C3O?NE788&:XR0TE[WFM3.NR?Rc@-g):QgXOc7B#K4@K+6+>FUCGSMX^aT,;
EQ_X(RTB.GY6IB].5T:>7>+-O5JUDG=-Y0D#b5Dc3G5^_+->YfN<;UHJ75WR65IP
B;c:&#MaK\:X9RYa6dHQ#7&=JJF_6]0Laf=&N@VD:6:aKD0>&VgM<Jb[]T5NNCQ4
DVO<]XSTE99a6(8?GI8(9f?Ea/#Q?J7D;&<)3QK/@B1IJa#gcf;PMTYRgJEf0VL(
U;(g(K4M,QA?.?9a\-O#]T3(31Vb+0f;dP=C)XQDg-4U_([Ke:611fb]^?T^S<H,
aNcVa#Y3E+ge;[^IWXT[CM?W;(X#?WC[FU@)J6//1XgY[K^L0NG+2#DW5>5f14:K
+_()=dEf.9a#RE\-&=fU\)TK=A:&.E8TdG+5HW8aQ6VE)&^&](\ZP+,)[KI/ZG,8
g>)J:UDF:HdE3(SG+8_)0&[49&3BHNg#]]\K\5M[_5ZRc;U9a<Q/[]H/SCgVMS4V
5gI3.5@?=PI(X35f6dIX&ZYA]1da53F8\#ODVOKcO>@0FcLcZL.0-7DI:UX.J76C
HB<D[^0_7X,U>c\0.2eG<2SUb>/,&LOf7:ef@4FUQ)\fP[IS3&=Z=Y/2.V64M@#>
KVRY[3c)f933A-W;g2J4(8FB:?,.,C;NGOaCJLWAc^cQQNWBR4]NX.)gV=&(b@=B
:)\d@+HNVMHSE:[#bc:LC3@fVff)..3&<D?WM\^N7JgFZBV#fGb7)7\=VW_)_O4A
:aEK]([RF&]e.ST)PAg6g(U?3=d=g1NAFeK#)88G[@<@F0HeW(YIR/N6965.Q)gX
._57_dA,D;3&0I,6=PT]W_2H_8[;J&GaA+:9ESU,W7_c&.QP9eD</E#T=MR(-)/@
aDb:Y]9Q@O#c2VMBMRP&?JS2DZ0J^Z?^ZBf4NV0d]NO?[&>#X^-4#(O(beWFAMKI
C5D7R()ANf<Q1I]7/4Q3c[/5V?.LfYc,W01A.ND#0JDIW0FZPF-G66#DEZM]7P+;
S+UBgfE60TSea#U69;YR9O&HL6UFH^eKe?IHVa7^aI+c21Z[ca198L)VW=8(J[G(
4];HX-a\&W,-dRS>gK##TSDNX9e2#Y\/U.F1W[,WL=OWN[2=V:gPJ10cC),IK&UL
SbfQ,S];F#_3;K<e;,9=NVA:E,@(;)_NE23D#GJ[PB6_8?f1BY3/JUeVWR)V,GG(
DAK:872\T8G9&Z^XTJ@NDP7J3Y9U@03H3dWgV=.OIP.eHTK_Y<g-V8dWNEc)6W-.
N7cG19bZC-J_c<CK40V1YdLfMb+5B;E,6YARH2FBd3BdgLN;P=NEcOWWGTA)RYK5
Sgf=(WA-BBFN&=T\<f[0P?5/W#U.W77eJH[.d6fD-V(+.^SPV8CeOW&1S?AS[65^
KObd2:G@)FD)=0@H:-F??9PT/T#?<)_O5e[.35EDTY3RC>^UI[;;_AcH2f-HO/UJ
[9e^3@a,P/\5f(cW&6[1Qf.8<cXQ6^<42RMRPHWC:-N(2JJX+c66ab?H6^18_?79
BC#KaXJLV#.^ZTDI2SIPR?/5VIF35[1/H-968B/BP2=J48SJ_2A;(LLT0CC_WT0P
NQ43?5^a0YaQ#)9&_XU#=_:4M6;\4@-T;D5BU-+,3Q5M==Ig\KD3_?(E6;Y>.X-)
TS[[+^JS;\>MZgb=MQaZL3M^HJH2R1V22QN83ReLF99JN^76)7>fSSEb2N78dDeX
)eG&g\WH#Adf7X+ZK,C#ENe8TZgP6472-]J5f30R6Q2]]4H4V38)_G:ELU0QcgNf
\=@Q62TBT[/)-D2F?b1.7^XJd>W@.]\(<QSa/d[5Z@2g+HD7BKFDU/^WGQ:KSH,U
P_R#de&e=V7S\aV&AN;IH0ZgUBJE?ALgV6eRb_B]BDWWWWKXPK3WO1Y=XQ+=dAOI
ZfL,208.J[\YLO2eb)-Eg1;+2U&U?SJWE8IcaI4#Q?0UEaG=?gGA4D:M69cS?OS:
FgLIZF(#Dd7Zc\MV_,_bf[BR)A1XF;=3^X\8Gf6FK?N_;?_#__H?;Rf;PJYID73a
@P+R-(d@=B&P7BTA&JPaO2P7_NVafd(-PLU,9N7]VM#/UD/52J:PNP5S9aZQYJSO
M2(G,[-WgDea^S)T9+e/9U=)UGXfU;PSWZ]00d?YPH8+S,daY5a=6+NJWQeC)=_P
c.ZZHa+CB0BQRY8F73+90G@V/K[&NA:_agb&.EeXZQRJ:Sa1.8AVZ=O,@dd\\XTc
D@3Q92A#c8V7a?0P8]dB-NA2Z4GebI:c;b<CD(c?Dc4N<2V>F68TZFS(-96F6Vb&
D&8Kd@WN]aV/C#eQ#Uf,S8]KZ3dJ+Ye..UKK/gQZ109WQ+>R[T_K.cS<AJII40cW
Z?,@bR9>,0gQ69TQV5f@0/V^M1LdeKS;2e&1bRgEA\MMYZ>,4GK?,J>TE^4SK2U4
BaF8g9],Yf\7GHHdWA<0?X8Y8Q(3aZN762#(NEGCL#PWJJL25#Bb;V^\E>LF?PKd
dDcQ.fNa7^81,T#[b3N]e<:V^##bbBaT4=BQ2^()L_R@f9P&g,ZB>e(4dX=6/_M6
86O0IVSJVMSUOKGTFS1TYa\HMX:3?X6H=7E/UW<I>ePVF8D1+5fR?4Ced]b@UJ(;
a?XYE,?O=QZI-Kd0JT.0?F5MNE&bO40]6Y?4Xb+L-7[JZ;DZL(fE7\MEPO?GK2)Q
:^1BFI/W2R^K^S&CT.dRLW<Td6W38?O1F(VD;B?_TIIfX6H=I7f8BW-4d7&D8?<P
@]YKT@^6P<A[ASdM-#Q//&W:&S1B4]71/_IIM.UM05e929L2IJ9@W+R[B>B+M-?U
DXe[aP/dSXF>E).X/_Mc9DKH:]S.3a.M257.8L)?PfgbDTA/NZD&ZEM-)DQgU.@2
]cM/U_d<6,<8)YB[[>BQX7Sb>;/7=B[2K^X3KfX,Gd6+.U<;&&F0(,#,1>,OL2\D
S2N6\U2R=>;Q+U5NKaUg;)2JVc-1@8T\MY=gcIfD+g[Pa:b.DZ^;.(@+3H;:RI,8
<SCBbD?3X6_IFgP/eY#?<2N4\CU/d6W)d,<3Lg_OE7V<,cUdM)d:\X+=cRTCT?6+
2H=8(+6FFTE7c/:c#d+cHfRO\VU1VV(?YY5G#WHE3@2[gTeG(g1<Y\cL;7_M8VIW
<[O6HW5YATUf^3(eeRDDg1MM^8b>:FcZJM^C;\QPGHPMK,\TN0Wg;.d1L83^X4Ud
Y7JS/SY+<&:#eb9Xc.U7g[,G41;<ZL#WUDb^]/PY^17/@:E5cH5@@aUe@VPc&)M1
cXMW<)]?bbE)&34-WJ&3c^VZd559YVOJ>SM7TQgE+(0,K[JJ]:_T=EM-5:L&0\&g
CV1fUX2dfFZWM4HB/B;SgfJ^J7-:#7N1eX^#55_D.N]H^K2OL7;-75Y^=aP<_7d^
(4E>+I&dQP#P_K1=J8UX5Y&P8JddLf]8XHc-M9-NMKKL6D_<7F4C+4Z_?US,8KEA
AB;-)>_MKK#]NYe)gYNXc2PTa/c8][1c&+\3,L75:(=<UK;JC3M[G+FIYKL6F(0&
,X;]c]M-(1:4D.RXEA?GOKKBG96eL(+-e,O@#,.1=W=4&a1BB_Z36V.4TfX=Ug[]
P^_45>H4ZCW?,76EMZ7(A1S=;>Ld#BXd2[1W#YBBA[?9[:KeDZ.N]ZSN5?dU1#D+
N<0\gV_(3=c&-4f&dD0PS>gM&;9HE>X:H\N?^R1(DLI4HX]21K:GJLd[Y>68K0-P
4-EfW9^N8B<73O\)\J14Y-KTTL/QAS-IfPBM=5=N=ffCGN(fDLg9HX(/>ZBLd85D
E=O;N?0#?dTR[eHcX+D-R>9DQRaS61\DJC1,N+,OJ]b\,I[Jg<^F9fH0:8>3gb4+
O=)2BLXYKC];1=5MF8db[c6XONK^ab-564J2Q+X5g^)-#7[259]9N6KdQgeQFF<2
>g.,d]6:?]/FGeTDTRVR8[++^bS-U0)A.6&2P[0>Cd:/__\]A8GW;YD)X2fH7C33
U0X9+Xc6+,?^2/M&CPM6ELKM;D).8IG2AQYB0#+4gB.;1H)Ja@S03c<HB.LBcW_>
GZ36_Lc-NfS4WOSCNW]Hg@9UD&CJPc?MVaAgX_IKV,1APSYYRN3faE7KdXYHX&NU
/#,37:Nb2E5b^RcB^,/>L^W.S@)(/<_/5&8&.4F_??WQ#TQ_d0f3S]X+Ta[BFD.f
2V&6Q)7U5?d/+g&KaXBUbZ5.+N7>9=8\^3+-1B2e@)02,bLJ^)547G:7E.#?<Uc1
XRFY&ee:\UX+:5cgI=^\^Z(BS5EOFG&aI#D93DQ.JR:,N\>MC6C:BN][(UX[9W@d
N<K?LA3aUTCGb4U87+2C,:8.A5C:++IO)7)-SE7;8e=&Ff?b.C6-)3aTK,[a\AD,
1.SBC1JV]TGbS.U9f/MAZ\U4UMLB,Cf-a-@YZ@Z5CF_96fO7(K#=L3JM^]4IN^=M
3fc[VN,J^b+DJ=g,.7D;1I&YDfO)VJKe_5OPde2@CQ>;#EWD4MW@c.OBgg(H#1M6
B;W56W_M+bW6]P3KS7I,N7W]5;8a#e871VL#2P77H(TKZVag6F+0J8WH3_6+_g;C
c]WZ7T+93AD@.QVGY)?^=DSSQF6UXZ7REU#KXT/@#ZA;M>=]7XCbAI^a_]FV=R>5
PKHN0db:/9Sf[HZOC:a58L](0a^-@?/#3@,9TT#7b0cNcROHN2CVY(B;e7-aB6V^
f8HM?Y18+4ETP^^-)-@[F88G:3=B)6H?XgbVOPT(-8:R)Ne7)OWU\6#Q<@,ZKWG3
&-03@Jc/B\R+d<0\O(9PE36HJGC18LMeRL8FfXIA__=0CT0NX:f;LRT3;9-QJON>
aI3UITTA4PfZ[.eJS]SCT=O\XXH[VTgI(7<7HXAHJF#)Yd[A>]a:4&S<[fWWb>gY
J7:QVSE1I7G^RO/E(,KLT(-Yc1TL?5d[J]#bES&@0Z)Y8QKT#Y3g=6WbNEY]M[0N
XG9VU=J^6<>&\F+M4T_2G&Aa2.^R\JJI;g[=CZBZeV2<-&L_A,^fV0fYB,6:fT&2
J,P)VZe)KEZb<-IT?X)XC]K#I\b32SOWS+O+=@b8eHH48A+1b)8BJZV_F+6bYRVS
)C/P@K]@V=fdJ)59D;cL,#KZ&dV.WUNU_<:++73_e\0;N4D@A3UbW\RJSgT5[=?2
;1&3TC@.01f4W4V&MY]&K=1TOM3a2@0PAS&MQ90J:W(&RZ=(Z2Q\JP7HG/YX7AB2
G2/0R:^40#0#PZR[a_SF&V:cG8:>1=CK:08D\5J\REf<g<Z5M@H<AHdgSG2M/)9A
PD[J5@B#)L+ZM.L?-?(be,>T@]_(bc+][\fIV1-R5JD>HJ7bf].9cNcXNJ@L?2>&
>3SZ1-#/K+7F;Rg0ZWU<Y+,_^]+E/2]>]MV+>&OV-TbR8/(5UWdEI]NH6ed1VAL8
aIbJ?[CQBTN(;eVC:df^>R6I&2/K]aA=],/MF_=F?[]F__9Eb#3I8[5UP;eF>a+C
06FJGCJgSgE0EPFBTGOQ>U[6c;5,65249@;O\[F2K<NcPAe;G7O?.b-eO,2JP[HT
d@\RB3J_FWFc5S=645WFWgf#MC-U&:<J?/B(UT)LB-=D716_=7UXeK)(8/P0XRaE
=;3&EU]4O2\@RV.]5>KIC/XW;MP^PH3H,X=K#E)(/+W=WL[1+S9+;+ID0^(3b<8V
SHc[U/YA[HVDR?Y0U0],+F.@2HB-SdE]EX(,T;A=Q)NC4YCee/W.b-YQ-_eJ<0Vb
/W#b<b6Ndc#;S=RQ(?3BPe&(D)NQ,#M,]4C+a+aM_21U=G#C9d[Ye+2]Fa>4+V1Y
?DKG-K45Q4d?8HdA8^8)_\;TM]DME^T8T\T]g(F>@c_73;.QMP-@-J((N4F#<B-5
dR)+4G_:c\dN+^A1a1[L,5&M-R,0&S\138b0,3?K=Aa()a/UR&#<#_d?c;VRUIEI
D?g@0AUJM0&YECCcS&CEMaW8D=,9WXPJ#^/CKG4=Q><ZQLbY;bMKB31fH^T(09#K
c76dL9WMBL6,F,.61=>8]8SGT3<7bGCQQ?18)bZa7R3ggac;=&MIP>+fa[NBAK:S
_c/.eVU=,fAKENSUBYc#?7W3Z_MB7HX-2^d4aFfC+I[RBFL=H3;H;9&WJaM#[5->
7)9&gf@0P@,/.0IU_NIA9HH<]J.aefDXd5JIf+R+CEG&DO^D@QV_abEG=.f#K^ZN
R,OaJ0\93;MFSE7909A+KZ<&;+A67eND-,4@d8JV,=EL1f[2:1\D.H1+/a/YO-E(
1,3dBAW4cTb.N8CgG@9,&6MK[c#g6b\5]:L#;0,D=@V:OU/@JCe+ZDM4@J8dEcaU
3&0G4EBdd3.4FF/9g.-ge)c,bdOH6O+:bfJg\\d@eZ@?.ARSJ@Sf@Pf@fYY]&\^-
83WNA2V1Y8ZIg-f6]+\V-L0HP+G#\eQ8fYJZ8bOc82Z/?8PVO^/A.>f)eGBK78@[
7^cLa8]R\LSd1caP2_b.A,<]LcZR30PHMYV,aa0g\fPVY@<&\,3#1.[]UO]]D+Fe
O;6<WPV]@EN(U\6K<X7gF2Pd8]E7,JK1EGBJ.^1=V2TTgRC3a[a^f][8],P@\L^G
KHc<=C=Ec3#?_B80ZbCE3B7D/F9;-ZP=]1gfM@gDB=de^E&80E#<^H<H.XY],bK_
0Sc2)gC\3cZc?9SUSU9?.=Z#+C&JGBUe3I?ag_X\;78defd<QL)]LG9GS@.T.PEe
5D_B.KDBDO,8HYT>SL0[LC>T=+D]fdS3=d+2a]2811NEX<Y)EB/([G#R^I(<#3Z]
17Ld^/G>23>YK#>(Q=_KN(D<e2WYeg=(=3V:+G@>941MZ=?>3)ONJFga#O(ZM3A2
42+gN6QE;,P-Y/YBLb[9=:R,P\=K;ae&OF+I>eT93K?T(#2S<EUU+XaE0@^JF78g
&Vf:_;A2T4WAagNf=J[E2+d+)9]df]PLNOgI19a-Jc&^XGYKQM9#:)4@dOMAF]WS
A/7K:RPD:BO3D9T6Y6.1?(d@g3DU8\[g:&#6)eOVXQUU-PZ=4BM..]UC6[Zc4\>f
aR1:<>/HXTT^ZT.eJ,5W):J>GFSM]Lc.0fCN]D=6d]0cP9^8fffHfYCb@=,#BK#g
IeR<c3J-BL:K]b_3KT/dPc;XV8A\3[fQ(/SS7E/5b=A^<,9[Y?DB+&>^b:@)2KI/
#R2;VX;EbH/;4OBIf5dd0V\8>2M#KU441Ge8V\F=Va#8V8C#+A_b\#g&\D,32M:7
M0YGRfV#a6I5/@@=BM9-KbU9(O=Z/]7/YScM?VCQ\ZeFcMe^-XS]NMCT]8NVHS+F
OKBWe9^Ee7-^-@d5_HKW+6KG(:A)Y=BIO;Wg55ObK_CKK12P=9MAY<4G(OQU1T&Q
=>>=K25>KaNI>2[J]ZZgA^;9If^LN472fG7)HOB-PUQLMUaNYKP9d&O#KEV7//5]
XM[#W7Pe01NZ.9fJbJW5QI-5b1-eeZFMFY5gMKC<H+O+R&KQ3T>d+)gQ1D?B6,a_
AR,W+&?X&TVd^KH@T+\c);;Dc^/-G:/5HG:)E79;K=EX.3aCV--_Jf9OW;D-XMc)
Ac0Z9d&9Z9<b<UE9fZ8V,Bf9Q4#]UR3Q7O4V>67E]@c5EH1;7YG#?:\-J#^ETd#a
P@E+O<I]WYIB.?910FW@X7W2R2:;,LO60GMEUbKLXRcLX\G@7=#SG;6KeCPX7Q@]
Xa&[Id5F>WVUf9W(<d(.<F8JM?.f?38MFS_?-S63(NLRgSP)3R\R,KgUgTg#:A,&
AA^R3](8>FL\AUVK,WS#,FJ,A.0<,(PF))?c,)R>EVdeV/,JbK4H8D)I1RaS:Sfd
;8,37>JUGIWR_E67#C6&4YSO=dDGNZGaTa/B0P5A>;400M:9PZ;gZ[VG\_>E(6cQ
H[MU/ZL/+cO_X-8,/cV_d?GXK</\-88Yb\KLCM,_9#Z/8Z)+gEVIg<W+<WOL1<:-
@WN)WfRcO6g@.17J<+S9MRR8N1TA=)M3W)OHQE[,6O&d]9a(HL;MYG9DMPe7:H/<
@VZT_9cg8A^77I53@BH+>BZJI4/1.ARL+AaDdBIJd135@6_:5CMZ7A5X/316\=N7
1;R^Y_Y3g_V3K7Wbg)4UC3MDg,;-NVNce:,/=@VFFCOGBX/CX^DCFU:0U^O]/fMF
/Y@>4]OX\(Q?FZMQL06H7;O4X]NFJ.?2+6F8RHg5>=bE9S^FZPdWK,&=12Z8A?K+
E0WX(U?(dDQ#L[8B/K9X0AKIDQ=OZ(>gbHY18LAM\=JaZe31b1&097\+WEUS;d4M
\de6^:_dX:6GZ#URE7BN..>8gK1;;81=\&.gec-OaUCWI63;HQ<&1M_[XSI&FdVS
];C4?K:@VfDR_A&f/I8Y#+dTX[<EVSX(M=^Z@/Q54B7T=Ab0?.K=G?aaH&eX0b,(
8#ACP,O-b5c@D&5]2A)R<c;e,4B+Z+]R+F1aWCT;X7Kg@=]VUNK3@Yg\2Vc23^MZ
/&O\9B9T/A1\C<D\&#R94(6:E(^H?C8@#ZZ&M&)UbBZ)D99#CKO<>XM&9X48CF64
:5HgV7A#U@PA/-bc<]Yb4>,V]d+CZ]dY2c?(&.ZYFZW9f8CX3R\[U3_a42G0_HWI
gH)2ga9c&-H[NY0<()^3ae-A1,Q<JTc/V<g[;SY4-H;A=93+TMU/X#2;A[J&f4K^
PDbKUXU0AL47,UN+A.HWD>ReYT^::]J\&F6:BU@OPTU;cf4,\O&)>:8IKBYd([(V
+?>IMSJ0XD-XW[L\QM^VL9GBUW]3Ka:fA:OEF@74fBGJB+g[ZGB(BQMJSL=AgPS#
SGXcL->ZMXGXLV/a,d^@R+d,F,f8HJ#PJV2gP=AN/f@+_XT\[(HEL^(4)H]M(,3[
^H@D@6F[&U<fU>daP4NGDHDRJJ9TQ^b/./TQ#B#N8J:c<AKJ,_2I;XDeVd0Q>HdT
,\#0ZYPNFH-gcVCg-PU4,./R\RR2]09gXG?d3M2b9aVFZRZ1UfY>?FgMc0GbC\BX
Sd.QF:92;=/?U9/IX9Q-9;M_K:ZBc1J5U0FZea]<)fQPFd34MUE9bF.K(]ALI_]2
?UZI[BAK5Oe\4^4LANM&e52X)5+(d4bWBBc:977g8cGZJNMJ[S;R;EY\QVDS]W>Y
(4e:8B78WKa[;6.W6Z[cbHS>?O<861FD>.M>>W3.@\I5+Bg2,):F_2?]aQcYd.F&
>4He>-3L=G)dQd]P4e[0ZSB_SORPaK2_eg;dZKML;>5Cd\]S0JdXfSKf,7;;@?fe
5PVg/#:+K^OILMDdJM/E7QPB?X];dZXWWX0\c2HgfgEB9V:T<TE+;,7JK#<+YFL=
#C[e=P)PLYLWG:+]\ZJ^?&W2aER9-2S=-_NGA/R^KUL1]O@Od4SZF@0fAMT;a#K0
V=H9>2(S:ZT-<ScgBL>&f=K>?aYTV@^D[KJ<.ZF]4V[5faC#d/IJEgaV(]8/<-RA
0B1Y9JIR>eX_J1-4^&Df>O/CQ1B?E\K8\=+GeCPVZALe7VCGfXO=&&L<Se#+BAWf
C5&8RC1A?d3?aLZ<K,[HIY#OGb:&/:_)ROJ>\M,9SeAOd:;/6dJGM9E>-#<3R]+\
b/,:Wf@MHf5eY_W670\)4]9Z,@g)ER5O8D=N_&#_Ufe>QgM<fb2J-ESH4e&I.6de
<5FQgg\LY=/S/fZef7ZVCc1)e6@8)e.=.&)5X3F0UHSE<F@6XF5JbI8O&/C1Y1-J
#U[X575a<d2IMH?=>TeSHTTN?eP[O<[4:g&c?F&C+e_#29X:dHHB7Rc>1DI5U<&\
9gc(<MCef3[f:2TQb8F#-[L:6_7YE)cEQ^1eOE:HI@BL/Z((gP@gX/:6Re2g\S+]
R6>&4BfSGQ@b4/H\MAG0F<6b7,ffIZ.(07@0HN@6F>RD92fGW.(gBE5M]Wd&&a^H
L@BCZeRcP^aSA^R/;I,3b(+D[X+_:9c4P=2S@/@8:dIG>.Q?;=4G;N>>>/CRG]HG
dP=D/U+@;2Z>UD<Bf2S^e\2AMQ47c;ZA1d&UJ64[13#eU&6&Rff@1gUJM4=3I7N0
5)1SI25<>(\-QT.4L/H/B]Pe^J]gXBF/DBBL?[5G.<4.>afYF75.U7?Zg.X8R5a@
7ARU&XAUX0Ic[-b#DdVZS0GZQI^&S?e.XL8;/>,N6?&,d@9Ra,#7X2XVE.+5>><&
B\@@B7gFR5[e@KRW1[e=8H_U-,;:eLg3D[G7N-C(97<\]VZTNd@)BT2:<&U#Kb>)
<cI4BK&4_,,9;O@?=7eC.RGUV>>8--LO<((15(RW)LCN#@:5@\\47#8<b]Ad8-#L
I._?G>d,\;PR(2PP\KN;DEXCRcdPE)5-_GGX2-A&B+4;P?2G-2a<=1\KgaJ<b<SW
(K#TF[,g,BL:_:b::1MFM.,,fg9#PT:+1O(3:FJY-V4+HJO,Ob2JL:dL7-8-cf>f
]NX8,OO,E[;>+HR<R.[Q+>,.3fX6#KCKegN\^TL0D)QGaG)D7d0-NKY63]B.UR6#
8?DANZYMB4M-]CVB2+\BQ\6J=cDQ<QLPCNV?(K2eVHL/5ZDQbW49)FC4K#ETNXg6
cd++I9JKTP^HX4B/H:5ZBaL25J^T<F>[WM\^>g?1+E[W>SGgV4CCbUC38L^WU8Y&
RP_(G4RMSQPBI)dRGITceJYSgbg^YgU+NGP=\b(-\1c5,;?2?H,:\+AG85-fNUMU
g:IBe:4Q_N.fd\-K]OBaXYV:Zd4U:.:QH4Y9Dca\<^4(ANOW,_5cbfDe9QPRI^8E
8Hd+D^A6GG\&R+WfKQJY@?](LQQN_Z1<0&V&Z>9f-RUF<L0Jd=cg2#e4E,6?73ae
cA)AV#/CRJ42?:NFM>AN[,U+M^@M@gP#Q=RBB5P-+[Sd1M6&;=\@aYI&#3J?FbgO
:SLE^O7UF(=[,?+YCJ=O7(fCA:CNOJ<T[Y2Q5OR9337@OGRRXc.I8_/c,#62N+E#
:KMa/d-1->G8W@7Wf->6/78[XMZWZ0AD#AG[7.EQ(=Y1)#_-X1:H0(4deERfG=0g
-8g;_:[<])O6fJ;DSMG@2Z]8EW)R4#TSK3KeBB]]bHCA8FMbNXNM/T0P,+B,ac<N
f:;T)35b8CPObdU+]],15&SbDd?9?4W&Z/]/Y_,6Z3P?MZ)OaZ^dZ/EMOY0d[/X[
g-HT00]2/5L:?EOb#1>-;Za0Ga)f>>;M)gb\.H^g2<0eZB27eI/N4SF1)KDEL2LL
Z[).S3S;4LJ-YMO\C?<QFP4+,Z;&83:3@>87(4JYZUS^MPK_^>JYUPBV1/b6^#?[
D-eDU8\XV^BMY[/(Q,Q^O\DX[ZB(TG/=gT(8Pd=gD>ce8\K_?KW-HR@=2GKd#fF^
-)8D8[DSaRB/J7-Y;20Fa=R>e#BSOfe\S81fe2AaDE--Y<T_G^7a#WAgXbK;+\+g
Y1)\=E21OQG2;e]ZZ<J+>JaBIH8LCC;(B@PR\WFT<SUITFfNPRZCcLABGZMR\J+_
.LaVgKgCaYbO]<CXYCJ#W]2:J<NX2HaBW0+B2Og&3O;#[#=N+^=90bb0HK9.\,S_
Ng1_>)>;UXD:8-4d/^LEOIW/75)Z53X;19UGM(#/89X<8#=3=d-UX4T+Y;&/PYRe
@C\[&]S8B^+(g0eQ6):[PV6XeGL6BA@.T59P,>JRAM\S=XQaebBLH>H^,(L6+B3Q
>Y^BG_2WVEabZ8<JV&L\7^_]U;0e5EeaRXg1>9+.DbN:1f-LTdP,:(AKe\P,3.I&
B9C[<[WOg406\-1645P\f90&&WOH0CC;(353a:4#7ZML:XI6)#<=(-7#F+F,]f_d
Eb4,^g)&)>IA>2G_^Te5)bX5Y,M4TY9=&]O2fP@Sa;S6IcegV@SgXT43&_G_Ad1H
-[(A_b,c<b(eR(7Fe#eUQE0BfA5&.&3;KH,gKGYe&YG@826+3:<gC[G]:gRQP3MS
d&][af_C5?64G7?&J.O28,IN1+:9\YKZYD.AJ9FG@1=@7(O03gZ]KM8#TK@.;<TA
^+3+dY]BNDAEG@GN@(M)0NWN.BWfT]Y)VdR7T=IgIKX;?ZG?7_eI815RA?D[MTTJ
KNC)3^IG_Ga_#2b#>@Y5&&>bW:>K4^C44VHAD<8gYGRP?]1BYW&ALML6/KP.+ZD^
\4I7UOd[,<8^5_A8-H-Z):7X5RRDYY^>-WfUVUc?M9RRMJYbJZ\@.3-7Y+aJW^XT
EDZA.^_C=R\d??Q/>QaDVeHbcWH[H+NM1K_\1g_->a[3/))^DQbO.6aMN<aQ0.f6
2QEQ,V[-N1a(d(QMS)TUOP=1aSg,;bG\O&\VeN0^U<@73CNa:FUL;EI5PVLBHU^8
G/=Ne8R8V1]T#>0U&eRZ977g]W7#[H^c,QEY<)X?.@-//D></Nc>deS_N#J4MS\&
GA0EfQ5?.DZDH_UI7dcKX\2DZPLDc/=g?+b:>JB.4X>L_Q=]B5;KA]G02W;5[8Sd
Eg:dL+7_R\;6I5g&^\H]MP6_g7S\Adg&Vg(1_=B9CNDGO^OT3e)a>-V-M=))GJIP
Y)1Z\V/AC_fGS.0<bS(;8,28=:OAW&_Z.b4?B5_-.dHJSbA-E:,F6C;5&W66@;M<
3_5^f4bS\(PV\aUc,,?bOB9]4GE>]02+DGf](2[UHVVAWQYABW=PVMM_Og<#NYHT
>E76&]bNS57)S5Q[;.Ld:]+BSG:=R-\[^[^_c:BPO-<UF31c6fN6V2U#O,A3&X+>
XcWNS4>J/I,VA34]ga.E/?#?0?C-&:1CJ?,NgK;3;#]aDL4.)QY^??63-MJ>7+.X
aU1ega[_6_Q0\[N-=.-KJFGf2I[P_()8_LB\8_^K]0DfT?9BN[Ag6)BUB3XT:VOZ
IJA\\a/c)&Ae+D<c5cJ2NK8;;XJ:OJ^ZG9HLQd+]OF1c?SYe^J9IEM(:C856&-aU
c?M\UgX\G0->ATdN1=^\[OREY\59=fNfCX1<aa?P7,MQC6Q>=2;VW^)@]11eU#>.
MKcJ_e4EJ@OV8f+^4GPPAM[&C:aaN.eYJT>PRSQ5ZZHUc,(2.R;#?WSd-/,I#,E#
=O8c,A@125FF=>-Bfa]MY+e\A(_;T<D2PIcC.2D]>SQC=:[^:9=eV\+[8J]FgGB-
C-7RWU[Ddf96T1D&c?Pf_TK8d]e4IVTL[:RB>@Q(4:;WGFA_MIRAb@14V\>9dN6(
C-.-7&.S3?D+ZF+@0<1>(F;X;]&VM.&]5,N#JNeaa?>\VeT]ERX-c#cAAW&6DW@0
W7)1IZ40<5]df(a:ZCf_Z(O5^)V.__[VIY\AD&FW7FW;>BM3XBR=Qf&KG3_c].:R
VYV.U1/7E=fG(^[Je;OY<g0P=QO3(#V]Zc;c@1LICdb>PDIfN+ES2X9NIfGfeZWE
P,=-RQ][C.=gO)/5E-OJC(_OK_Q.VdY58ZC\a4A[YM2)((8<g;C]bK.@C#6L4D_W
#^&]/IOCIeQST^::8bg\f[Z\+ZOINc^MT_d8I)OD1gX75X,^PE2HB_BeUC5X0\F;
&aT,OYWE#Z5ac\fe5b,A>>F/f:)&K=SE/ObIZ.C9HYcN55-]XH-SFVD^H\,Dd5:L
6fT#:g0+[5g+#7C=BX81cR?HSJJ._LdN80[Z4WFRH1:O:D>d7;Z7^4f(+,4cQ<@_
AC>UQ3D5aKV2R<I#GccJ8(V7Vb5IHS5/XY?Y>V0IG>V&U(A[]QGECYC5,4?]1^),
a55T7G+bNHgCK1+]E/?[>AZQbH5f1I,G@[/4aXR<DNICffAFD\CW1;1/Zb_SQ:T\
?aT?>\a48O,Y=/FGVPG(TgRBDP+#]1V(JW@K(N7A;(Z#RbXGZ;=K=G-Y_^0&&HXL
Pc#@MZ0J>.JD)3Y,0fSbZ\B<=D8>VDC<+ZL^GeCbN+6L>=)QeJ?4U<MN;JY(eZP=
&IDSW6514Z3gAR0Zg<@TUS&95+cUfP[LIIb_]/A7HS@2YK)W,e)W0WY;#gGN^fJ5
R3.\=I<O.9f+:FVB.A);TEC<,Ff&g@[DQW#-/5&UFXTDcACeXWN^[INA/];5:-+/
(OdXG/6]()<17<3dQ<6\.?]^JP;MSJ#IF#X3f3=G2DJM^_>a)PJ/58DX=/.#aWA.
7AI&TYCX<N;,M]eE/;Y(3LB5]e4E5\H/4^@.K(6FV_H9.G\S6IY86f[^OH.@F=]N
]C\=C]8SLV;M\f4_M0L0JSMUZ+HHN1@\TL&CI4Sc-g\gL4=L;&e=J-Mg;]\/2fJZ
g8(gV6+P/Ke<Y/]LOPX\?XX?BG3(&K\ZN8B95T0UJA3:EdMD,b09PY:&-D&5R>?Y
N(?L_8P2DafC@R:RNe?7F+2@2aX(6eIVJBB49OaN,;PC+19Dd^[e2,HTPa];:9A&
T#,d-:5G7bH)GAe=ED9H99NP/5]c--M?@H\6G;_AW9K;\,F:4U;e6&:Bg\g,^eg&
@QFWG:D.,_UaBWDJ77^[e2B@]H2\;+W=8;>V;N-=/:K[,B\_6;cIOgU7.>+O>QYU
U-E-DTR(@#LI:.2^RIF<@]HR)AAd5@GDK=&?2d,A3X[9WgD,[0FK_eX-C850_^KF
:fY>,O\bFN^Ee>IGV:?ZEU&)VDS9#B9ZO;L8f\Q#\Z^BSN;/)F^Y0(C?H19,aN6C
WW>E@cU8,QEX>_8X>;\.>BD<P+GFF@UK\_^dCaH,:8,fQI5(S=JLC-<49,gH7Wbg
T+[]MA=(W]_a_R<^>Z:2^_@^gR12Vf5aP>cY</]PH0\cg5Qf?HE=>,Y\_NFKMFA4
WSO&[IHAI=Q2\9Gd@:K.@V?G5C?aT7.A2D]f2;UZ(TU2F#YS&:.becGBBD0^.H]g
023/6>db>LFPSPDUQ:bDD&[2WagI[Ba3_g:^+^g68_GIL8\<@Fa6=U[=dVLNC3M2
],J_L20_ZT(f?,eWeMFW.S0AX?Fc31;bKZ[Y8=Y#+14+<MUOJB1T=VSg)g=ZJf^&
Z:f&KM)TF.3MAVSW/D@X.acPa/R;3#;eCWCY+F\,D[[U0HIYVYR1&>9XE&L.,7&N
279N;(E#?^(bCM&#1O8,+&MTVa@;,8M0T(\E@@)(..9,T#a17@[I^X[37GP+?>V1
>PD4[[Y/6I6M6<CTgJNfg/2#ZR@(Tc\cG_6(e[08ecQFb_aG2bMSRU+Q=8[=:7VA
\M&WJfU[=&2I]W=6U<E389K69+;UM-9g+T:],_9IZMUUDY8-,NW<45D3A^ITEDO3
3H]fBT1(_E\:bXKXN4A[)_e5A1;KY@_1<E7@8aFXWQ<+MM)R8^91O32eacPb1@9T
a&)X\W])._9eG&g4)d7PIT/#Y;OV@bCgE@C9C1QKCB[9O350\@&^5.6,7Ef(GS62
-4=aa:B3;_D4E-b,]:eWTRYAbPTZffQ6=S?_0aGZ/LW7fPRVFGBBEDOg7@/Z-&IE
HF2Ug2Aab<AUafa;X22f.9U&362)PLO5J;5^DaJe8GZA,&f8,9U=?)Jb/P]3\b]5
PWF1X+::9ONO;g;&A<UbDNMJ1/(JD:4UJVC48a@J=cHD]=(#1.WT.I0AFL[dFKO_
GS7<fUW/BCB-VMC)PI73EgT,^2?,GPCCJ7,0dIMdC_T8_ND3Wa7/[51gIV500(0c
6AD@ffcCbO(27TfOPaN8;+b])U,fX3V5C]IfR^.Q\;<&JaB(d6Z\=G&0bb3JVTXQ
43@e5\g<WD6Q-FAe6H@@AYY^EH)EFNYN;Q6)E+6?LNCXZ><Y@J^Z<<8f=_Z7a[Z;
^a8Eb\-[-=</dTG9#cgI+-UQ>c5(K.D@6SZO]D//2Z36LQKd7TF3JDBK7R<I+@>6
AEbVYE9e7@X>Y:=DJG+RfHQ=4>1G9gUGHUK4Vf77Y)X?KXB=S3O6g.)fVfZ,GIdT
b\TC6/W)MV,f:&@T?SZ<<1?aPR)Z3<K@2O+P8B=;[)c,P9(Tf34g@;\3f:^a3N,=
+L>7(Jc,?<#5-3?/5^1RCgG7M<U=16OZ.)TC\LEJ^L+c<@5^ES)UYCEXEFQ?81+1
27WO))++_R(J=S;>P-VZKCE3[EK8c84@]QY>PD><g#:<F?24fX9-33P0+5L+(W8W
W./EDf.N4MA>_81_2YN/8+gFV[B6dRW2\G3]cIfKIL3-d7/_HDJ82KBC2.<LO_AR
>F8LYb3K(?AW;=dL#Heb)IcQ8;]EM6<Y56]ZAM6L[&FIP)a#aUB=G/B0TCBd9A9J
E)LQVC\^.&Hg7fVP=bGS1e)d7/+4Z.G5NOEb,a-6e/2=H.;0W@Kb)RMV.cIY<g\-
47gUDcG#[f#M#5gKRW[/@R/cFF]0=bJ7>UL(BNK&1N66c;GIT_&G,6#;#+#=W0+R
ABER+\Z@fbgF6NFESg07^G4c)PC/@,[G3gGY&&T>56#1KHO#D@0K&UFdHdX8;)/7
PSQV.3b+?5EFR:/#(ORHS,S\DEX)9[>JZ13#].&5N6C1B9L[6+R96&?UMdLXP8cW
:#).T2MK12eG.\5@)c-[HX_,]Y:T96BQ;#61cR:VT6eAB=&U4T49N@+a(.N4,a+G
Ue7#1Kb4e[(K7R]NI03f;WP]\/8,/+BNL7CMdNLNLC,a/4@R>G-K;/6</T8ACNf<
#VLd1NHJa6e3JYSW,/Ua\?9=]K[aB1)7OaF#FY6HVfXW.#?0@CSP?0I@cHCMd+Ed
O.fdSBOeE)Tg<V(/23KR?BdT[?>RbOJ@Cb/W[/;+\=Y1R?/-DM_]Z4a_[b?Z=.\d
21RJ[fHS6J4\fK9TN@=TLK8B/F#da<b(.e-?OE)]_RK#JET&-+9>29,8QUYAI/X]
_.T_,H(_/d:7P8F=_fPDP6,OcD@V0+?0X:1)>FN[FXL(/,a[G;E6Q\+XJWF\#/8W
:GE_D=E5>HT5TA9:[@b,@MV\P\DX;_#f3Z1>JTW0<bY:RY6#4LB.-NaNa(.U0S2=
dJPR)_1T?R>fb&HK:BGVV9H)P>>3gZS#1J5IdIY86LaMI>4(gGA-<8dV>6SDbZU/
e6QOKJDfR(Z_EcF>H4e#G-IXA7QW^N64;_9ETXV)7Y-NR[G_.A)IZCN_Q[4V-3?d
41/>b1H5();E<^8#(6R(XaU1c9_RfE8F(E>g;&NdOL4a-K&LP5<?G_[>##DZ2B\?
G>[G5Ne48d0J9#3_/)7d91D0T5bPLR_YW-eX-Y;3gT#2YS)YR1cgd:TBO;(cR[2.
&_,A(d=B.P?ZH.L,=@ZbeJ20O&=)YMEXDA(9(JGS5:,gG^A,3d;.e_ZYY3,+]Nc?
\PP?b5TOJ0VeK<KR5(O@TcH.abf0,]?c1c?D.SGVOR<gW.PdK4:HB)Q/-g:A<E^)
2@].R7;b:RC1U\_OA1:cM@-/1gF5+2SDd3_4;?Q(e/\(dfP9TYU+6UH@8@H(&342
,-9b-RLIg5G1\WF0&\/H&Y)eHRO\1XMB+CY(SZ7\;RE0@W4.+?eAPOHR=gEK@AI+
-A0+-8_RD+RJNf+?g2a0LXS@dD;3dYfG3/^8QAcKdeJI\2M41e(?,QCXCO^JY?4B
G;X\=UH5T?GE9SF/_./]]Z0;NQe4-E+20,WVDM00I/[eM8XdfBN9f\8SK9[>Q-9X
fGb,d;:fdH+@>+>0EJI-Wfb/@,M0X?#/,[\E:JY<S&LS6S2VVMA:cV\)E&E>O-bJ
8;?Ue32dFAdaE<dd]fWXR_LA-PcID9U)A=C#N9g]UVeP0gJJ[Ld/=e0Ug82P9YaD
b,15Cf@]3TbW&I7W49><EINPY[gBD=C/,V+PHdM;WS1N-NRZ5P-;Z[)>Q3GEZ1TD
8:UFTY1A8f/)2eZ7\a-]RSW29C@I@-2MB-=g3+AF,K;Z<-<,2&X3dOG2;X;]AE0)
CX)0:@ZOENC-H_W7#?J._RHQX-cEWbZ;NYU,L3bg=^_BeN+J8]ZSRT2-2/RV5>N[
=V,_ERRXXT(WM1=eSU/<E[K[=L#Y?BZL<eO2cR5?WW0>:[NK?aVb19QN]8N7(9Z7
X6Y&K8-d_V,CL,O.;0ZC-N&JW;BA+;PPBOFdCYK0)f<PXFE=f\LQLVE6O4UL(3D@
E_D^=+\7;dUVK5)B-L+<bD-/3cZFaI]6;KKM0QcR/fDT@\DBU-IUg<U]5KTI[U#O
N]=.J?E+ACK+U1;HaDcRFR,61S,OZd?<.+(c?&&d1&9;\GNCX]Tc=AV]ID]g5=4c
2Z;Ac?eY_RR0dgQK>1gaY3cb6;-P0.TPa+OELG&BW,Y(0Zc\AgGR1NQ6I,=1K8ZI
Q,B#04VI_TN:]]4&T09J7Pa<\YD#K22MGefb\G:g_:L,2ZTI@0VXLB^4Z9#MV8R<
1?QBa+C6YaW,7/dO/P8M3c);[cGX8X01P:KR5J;T?8UW7L9@\JDDS1^Q<J?Gg>DN
>PN-fB]WQb05A<\Z(0c#.9E3X4Oe]Pg-LVG5=6R+0RWM<X\gBH.&ZB#c12:\c=UD
)V,R0CID+4c#HB5G(;NM9W>K.eB90T_#UO5b^@NPG+deCa&.VcA=]QX&WD[&,FSe
(3DgFAbUg<Z6fJb5ePB#bR2dBH.TRLQ&&HZ0g,FU:P8@J/DZRg0>fA69dWC<P1Vf
+Z,R:G<U/4aEE<ZTJD=V;_O>Q1(UI:7,@H#1+P->H>I4\M70]6D@0.cN:7-]A(6D
@XVD6B=JH[C3N1<@X.O-9?C)V8DFHEHY7B,e-,R8\e,B=4UX55&>&E1(L9Z:U,LU
2;TEf,^#N)58#4_=U2FM3V+0JZPX7@>QR@5BGUFfQZ\T,6S8W/T5=B0JVLO(dg98
_UX^8K-g,c\_T,fd7)8P+UMTZ\>fIL)a446fC0D[MT3aZ[Ze)RD>+A92.[IKLLAa
2G=PAdcG6^fac:&dP&@;&_F?^38;5.BAA_(?\cTXW3J&f5:)gIP-8HGP5I[cUC-P
BI;J(DQe_N5E_Ad-;BH(._.VP[]c(TJP]1gN>2+N7]6N_MPba5^SJV#aaEB^X=dW
-PH\6KN\PKAM\<^?1F_NV:OaSSC/B3>BCb(LZBb807c\FF)T;>M9RPSdG+A4@@>d
;Z)S::+]S1_Mbe5db>?GTL+7e0cXHTOSTJ,SEP3_(CTJ(RgLS6O,Z3Y4/?1B3fL\
AdN[+O10GLDR?OW<>dY6OU9SM,\VEdcP,-JeQ/b7f=7?P+T^A6ZNg_^cXdS5HJa.
gcb+7^A&.=(]\YWQ/e]&GK3dU\N(K.@g@:0Q8&JT)P^d-PFF6e)LR-4F>TaFT@:A
(&IS,#:3X,JX=b^+0-AbgIB2^HbESI[ZXZ2(I>f@dHXH,LNFAB@-eQ:/a3d5J_[1
2GEFFPf]ZOE/F;0RcHQ97+eQFQHJCWDgYCSIYM<AHZZFE<g,Z.0RHL5SRR+.L2EY
]8X)>Y6gAZD:KDK-ZMd\^.a,:&J&J^+&#57b5f;\P(C2\#[FOZ85D_U=_HfO:gSe
PA=[;c<cGgCNfU530=T1:922._8M37Z#)04V\e[W_5BE9<T31XGL/>?GP,E?G;fZ
PJ^8B&8Hd:aI,XL4?KfFCK#/#0fd))ePT4LKceeIDN]X&.fSX(/5JUAX-7SYD#Rb
gSJeNI;]dB?F/Lb0/T0_[\WU(PTM5Bf\b8<&H<H.\Z=VRY)<e3ZLZ@(aU3YM)HTY
;?+^P5AR-J;9K1<CeWX;;d:+d?eRccRC3a6AP<6eSa8g@(SESY1T\dF(CQ?T?I.)
(+YE_4EOf,G:I9:H4YV-56=Q)bP:BIW&5d,H.YKC9:?^(191VH4_JNg[\eUE054L
&(e#-a&Ka=_>aM8@CSER7T=7:ADYKC?O/5XYN(&2E,OOC,4g)P=Z_4OE2S6CHS\;
a^5-9#2JCK0c&3a/6UEcQ73<HH<IS8\6AZ4BXMOP2^O#/WgEO0KdaU#4d/3+7P8C
SZ?g91GR6FIU#Y(>be20>8Q,BH:]McIM.Mb^N,cA,7,1P^;]]LaM=2&Q9ddbLgeg
gIaPe@>;M>-98;aV/IIGb>Q6GK;+PU<I^C>#/:@K_OBA#NYHL)T,ZDE?X?X?F/_C
:+gI>a?Q=3YJDgH)+D\W53QL[(6P1E-60<^fJ459f2FGB77>+a=Y(42<b+01cY>8
F8#?TeE7.6]4QQK+K6+d(be8X0ZfLIM^NC.N+/=c:FDKMF30]>AO)^3>:+I3IP+1
8EC@#Kf[&X_-]T+TGH?JeY.aZS8D;cZM<SG/f)@5GA\TMJTVX+5FDT,#Z=B<8,.8
eG&/9H]0/EB1/A=8.SX.YHL#G=7#9<WQUPJD6<EQ;V@abW<[Q>c#2A1US1D([[G2
IUdBd\).]2^3=&DbfQ/N6gYI=UZfJceYE=&[NcTSa3-HZD-5@.+R;[M6C8;O^Cf0
(/VP;I4.-;Cg\\dCY-++@P6XOTO/ce1WZCZC9+GPdeVKZB,<eU5\\:FcXgbYTGPe
TLMC9]<@]KP5+cA@Cd,TE^?ER/JJUJ-UCLG=C3=/J1JY5K6/ZXbc2cFBO==+bg_NT$
`endprotected
