module Program(input clk, INF.Program_inf inf);
import usertype::*;


endmodule
